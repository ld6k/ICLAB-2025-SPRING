/**************************************************************************/
// Copyright (c) 2025, OASIS Lab
// MODULE: PATTERN
// FILE NAME: PATTERN.v
// VERSRION: 1.0
// DATE: 2025/02/26
// AUTHOR: Yu-Hao Cheng, NYCU IEE
// DESCRIPTION: ICLAB 2025 Spring / LAB3 / STA
// MODIFICATION HISTORY:
// Date                 Description
// 
/**************************************************************************/

`ifdef RTL
    `define CYCLE_TIME 40
`endif
`ifdef GATE
    `define CYCLE_TIME 40
`endif

module PATTERN(
	//OUTPUT
	rst_n,
	clk,
	in_valid,
	delay,
	source,
	destination,
	//INPUT
	out_valid,
	worst_delay,
	path
);

//---------------------------------------------------------------------
//   PORT DECLARATION          
//---------------------------------------------------------------------
output reg			rst_n, clk, in_valid;
output reg	[3:0]	delay;
output reg	[3:0]	source;
output reg	[3:0]	destination;

input				out_valid;
input		[7:0]	worst_delay;
input		[3:0]	path;

//---------------------------------------------------------------------
//   PARAMETER & INTEGER DECLARATION
//---------------------------------------------------------------------
real CYCLE = `CYCLE_TIME;
integer       total_latency;
integer       total_pattern_num;
integer       pattern_count;
integer       file;
integer       r;
integer       SEED = 82;
integer 	 num_patterns;
integer 	 pat_id;
reg [8*8-1:0] str_buf;

integer get_ans_i, get_ans_j, get_ans_k, get_ans_l;
integer mn_i, mn_j, mn_k, mn_l;

integer res_mat_i, res_mat_j;

integer get_cost_i, get_cost_j;

reg [3:0] src_val;
reg [3:0] des_val;

//---------------------------------------------------------------------
//   REG & WIRE DECLARATION
//---------------------------------------------------------------------
reg [3:0] delay_pat    [0:15];
integer   edge_pat     [0:15][0:15];

reg [3:0] out_q_source [0:31];
reg [3:0] out_q_destin [0:31];

reg [7:0] ans_worst_delay;
reg [3:0] ans_path [0:512];
integer   ans_path_cnt;
integer   wait_out_valid_time;
reg reset_done;
integer best_cost;
reg out_val_ok;

reg     visited      [0:15];        // Visited flag for each node.
integer current_path [0:15]; // Current path storage.

//---------------------------------------------------------------------
//  CLOCK
//---------------------------------------------------------------------
initial begin
    clk = 0;
    forever #(CYCLE/2) clk = ~clk;
end

always @(negedge clk) begin
	if (out_valid === 1'b1 && in_valid === 1'b1) begin
		$display("                    SPEC-5 FAIL                   ");
		// The input signal should be zero when out_valid is high.
		// display_fail;
		$finish;
	end
end

//---------------------------------------------------------------------
//  SIMULATION
//---------------------------------------------------------------------
initial begin
    file = $fopen("../00_TESTBED/input.txt", "r");
    if (file == 0) begin
        $display("[DEBUG]: ERROR: Could not open input.txt");
        $finish;
    end
    
    r = $fscanf(file, "%d", num_patterns);
    $display("[DEBUG]: Total patterns: %0d", num_patterns);
    rst_n = 1;
	in_valid = 0;
	pat_id = -1;
	out_val_ok = 0;
	total_latency = 0;

	force clk = 0;
	check_reset;
    for (mn_i = 0; mn_i < num_patterns; mn_i = mn_i + 1) begin
        r = $fscanf(file, "%d", pat_id);
        // $display("[DEBUG]: Processing Pattern %0d", pat_id);
        gen_delay;
		reset_edge_pat;
        for (mn_j = 0; mn_j < 32; mn_j = mn_j + 1) begin
            r       = $fscanf(file, "%d", src_val);
            r       = $fscanf(file, "%d", des_val);
			// $display("[DEBUG]: Got src:%0d, dest: %0d", src_val, des_val);
			out_q_source[mn_j] = src_val;
			out_q_destin[mn_j] = des_val;
			
			edge_pat[src_val][des_val] = delay_pat[des_val];
        end
		@(negedge clk);
		in_valid = 1;

		for (mn_j = 0; mn_j < 32; mn_j = mn_j + 1) begin
			if (mn_j < 16) begin
				delay = delay_pat[mn_j];
			end
			else begin
				delay = 'x;
			end
			source      = out_q_source[mn_j];
			destination = out_q_destin[mn_j];
			@(negedge clk);
		end
		delay       = 'x;
		source      = 'x;
		destination = 'x;
		in_valid    = 1'b0;
		get_cost;
		wait_get_ans;
		// verif_ans;
		@(negedge clk);
    end
    
	$display("Congratulations");
    $display("Simulation finished at time %0d", total_latency);
    $fclose(file);
    $finish;
end

always @(negedge clk) begin
	if (out_valid === 1'b0) begin
		if((worst_delay !== 4'd0) || (path !== 4'd0)) begin
        	$display("                    SPEC-6 FAIL                   ");
			// display_fail;
			// The worst_delay and path signal should be zero when out_valid is low.
        	$finish;
    	end
	end
end

always @(negedge clk) begin
	if (out_val_ok === 0 || pat_id === -1) begin
		if((out_valid === 1)) begin
			$display("                    SPEC-5 FAIL                   ");
			// display_fail;
			// The input signal should be zero when out_valid is high.
			$finish;
		end
	end
end
// $display("                    SPEC-4 FAIL                   ");
// $display("                    SPEC-5 FAIL                   ");
// $display("                    SPEC-6 FAIL                   ");
// $display("                    SPEC-7 FAIL                   ");
// $display("                    SPEC-8 FAIL                   ");
// $display("                    SPEC-9 FAIL                   ");

task gen_delay; begin
		for (get_ans_i = 0; get_ans_i < 16; get_ans_i = get_ans_i + 1) begin
			if (pat_id === 0) begin
				delay_pat[get_ans_i] = $random(SEED);
			end
			else if (pat_id === 1) begin
				delay_pat[get_ans_i] = 0;
			end
			else if (pat_id === 4) begin
				delay_pat[get_ans_i] = 15;
			end
			else if (pat_id === 5) begin
				delay_pat[get_ans_i] = 15;
			end
			else begin
				delay_pat[get_ans_i] = $random(SEED);
			end
		end
		for (get_ans_i = 0; get_ans_i < 16; get_ans_i = get_ans_i + 1) begin
			// $display("[DEBUG]: delay_pat[%0d] = %0d", get_ans_i, delay_pat[get_ans_i]);
		end
	end
endtask

task check_reset; begin 
	// $display("[DEBUG]: Checking reset");
	#(CYCLE);
	rst_n = 0;
	#(100);
    if((out_valid !== 0) || (worst_delay !== 0) || (path !== 0)) begin
        $display("                    SPEC-4 FAIL                   ");
		// display_fail;
		// All output signals should be reset after the reset signal is asserted.
        $finish;
    end
    
	rst_n = 1;
	#(CYCLE); release clk;
    end 
endtask

integer computed_cost;
integer prev_node;
task wait_get_ans; begin
		wait_out_valid_time = 0;
		ans_worst_delay = 0;
		out_val_ok = 1;
		computed_cost = delay_pat[0];
		while(out_valid !== 1'b1) begin
			wait_out_valid_time = wait_out_valid_time + 1;
			if (wait_out_valid_time === 1000) begin
				$display("                    SPEC-7 FAIL                   ");
				// The execution latency is limited in 1000 cycles.
				// display_fail;
				$finish;
			end
			@(negedge clk);
		end
		total_latency = total_latency + wait_out_valid_time;

		ans_path_cnt = 0;
		while(1) begin
			if (out_valid === 1'b0) begin
				break;
			end
			else if (ans_path_cnt === 0) begin
				prev_node = path;
				// $display("[DEBUG]: Worst delay: %0d, best_cost", worst_delay, best_cost);
				if (worst_delay === 'x || worst_delay !== best_cost[7:0]) begin
					$display("                    SPEC-8 FAIL                   ");
					$display("Failed %0d: Worst delay: %0d, best_cost: %0d", pat_id, worst_delay, best_cost);
					// The worst_delay signal should be correct when out_valid is high for first cycle. Otherwise, must be reset to 0.
					// display_fail;
					$finish;
				end
				if (path !== 0) begin
					$display("                    SPEC-9 FAIL                   ");
					$display("Failed %0d: Worst delay: %0d, best_cost: %0d", pat_id, worst_delay, best_cost);
					// The path traversal by path signal should be one of the critical paths when out_valid is high.
					// display_fail;
					$finish;
				end
			end
			else begin
				if (worst_delay !== 8'd0) begin
					$display("                    SPEC-8 FAIL                   ");
					// The worst_delay signal should be correct when out_valid is high for first cycle. Otherwise, must be reset to 0.
					// display_fail;
					$finish;
				end
				if (edge_pat[prev_node][path] === -1 || path === 0 || path === 'x) begin
					$display("                    SPEC-9 FAIL                   ");
					$display("Failed %0d: Worst delay: %0d, best_cost: %0d", pat_id, worst_delay, best_cost);
					// The path traversal by path signal should be one of the critical paths when out_valid is high.
					// display_fail;
					$finish;
				end
				computed_cost = computed_cost + edge_pat[prev_node][path];
				prev_node = path;
			end
			ans_path_cnt = ans_path_cnt + 1;
			@(negedge clk);
		end
		if (computed_cost !== best_cost) begin
			$display("                    SPEC-9 FAIL                   ");
			$display("Failed %0d: Worst delay: %0d, best_cost: %0d", pat_id, worst_delay, best_cost);
			// The path traversal by path signal should be one of the critical paths when out_valid is high.
			// display_fail;
			$finish;
		end
		out_val_ok = 0;
	end
endtask

function automatic integer non_recursive_dfs;
	integer best_val;
	integer sp;
	integer i;

	integer stack_node[0:15];
	integer stack_cost[0:15];
	integer stack_child[0:15];
	reg visited[0:15];
	integer current, cost, child_idx;
	begin
  		best_val = -87;
  		sp = 1;

  		for (i = 0; i < 16; i = i + 1) begin
  		  	visited[i] = 0;
			stack_node[i] = 0;
			stack_cost[i] = 0;
			stack_child[i] = 0;
		end


  		while (sp > 0) begin
  		  	current   = stack_node[sp-1];
  		  	cost      = stack_cost[sp-1];
  		  	child_idx = stack_child[sp-1];
  		  	if (current == 1) begin
  		  	  	if (cost > best_val) begin
  		  	    	best_val = cost;
				end
  		  	  	sp = sp - 1;
  		  	  	visited[1] = 0;
  		  	end
  		  	else begin
  		  	  	while ((child_idx < 16) && (visited[child_idx] || (edge_pat[current][child_idx] == -1))) begin
  		  	    	child_idx = child_idx + 1;
				end
  		  	  	if (child_idx < 16) begin
  		  	    	stack_child[sp-1] = child_idx + 1;
  		  	    	stack_node[sp]  = child_idx;
  		  	    	stack_cost[sp]  = cost + edge_pat[current][child_idx];
  		  	    	stack_child[sp] = 0;
  		  	    	visited[child_idx] = 1;
  		  	    	sp = sp + 1;
  		  	  	end
  		  	  	else begin
  		  	    	sp = sp - 1;
  		  	    	visited[current] = 0;
  		  	  	end
  		  	end
  		end
  		non_recursive_dfs = best_val;
	end
endfunction

task get_cost; begin
    	best_cost = non_recursive_dfs() + delay_pat[0];
		// $display("[DEBUG]: Best cost: %d", best_cost);
	end
endtask

task reset_edge_pat; begin
		for (res_mat_i = 0; res_mat_i < 16; res_mat_i = res_mat_i + 1) begin
			for (res_mat_j = 0; res_mat_j < 16; res_mat_j = res_mat_j + 1) begin
				edge_pat[res_mat_i][res_mat_j] = -1;
			end
		end
	end
endtask





















task display_fail; begin
	$display("[38;2;151;132;151m@[0m[38;2;143;121;140m@[0m[38;2;142;117;136m@[0m[38;2;142;117;136m@[0m[38;2;142;117;136m@[0m[38;2;136;114;132m@[0m[38;2;141;121;138m@[0m[38;2;142;118;137m@[0m[38;2;141;117;136m@[0m[38;2;103;88;110m9[0m[38;2;119;96;115mB[0m[38;2;143;118;136m@[0m[38;2;141;116;135m@[0m[38;2;142;117;136m@[0m[38;2;150;129;144m@[0m[38;2;144;123;141m@[0m[38;2;143;118;136m@[0m[38;2;124;105;128m&[0m[38;2;78;61;90mG[0m[38;2;87;67;86mS[0m[38;2;109;93;111mB[0m[38;2;97;77;97m#[0m[38;2;138;119;132m@[0m[38;2;149;129;146m@[0m[38;2;144;120;138m@[0m[38;2;141;116;135m@[0m[38;2;140;115;134m@[0m[38;2;140;115;134m@[0m[38;2;140;118;134m@[0m[38;2;129;110;129m&[0m[38;2;108;87;106m9[0m[38;2;138;115;132m@[0m[38;2;140;115;134m@[0m[38;2;143;120;138m@[0m[38;2;138;116;133m@[0m[38;2;138;114;133m@[0m[38;2;139;114;132m@[0m[38;2;132;113;131m&[0m[38;2;92;78;100m#[0m[38;2;70;53;80mH[0m[38;2;77;56;84mG[0m[38;2;83;62;86mG[0m[38;2;124;100;116m&[0m[38;2;105;86;109m9[0m[38;2;71;53;80mH[0m[38;2;93;70;101m#[0m[38;2;105;83;121mB[0m[38;2;101;81;121mB[0m[38;2;128;112;141m@[0m[38;2;159;149;171m@[0m[38;2;129;118;140m@[0m[38;2;106;86;105m9[0m[38;2;131;106;125m&[0m[38;2;103;85;105m9[0m[38;2;72;55;80mH[0m[38;2;92;70;103m#[0m[38;2;105;85;118mB[0m[38;2;139;126;152m@[0m[38;2;152;144;164m@[0m[38;2;149;141;163m@[0m[38;2;126;112;132m&[0m[38;2;120;100;121m&[0m[38;2;103;86;121mB[0m[38;2;134;123;151m@[0m[38;2;147;140;163m@[0m[38;2;145;137;161m@[0m[38;2;145;137;161m@[0m[38;2;144;136;160m@[0m[38;2;139;131;155m@[0m[38;2;141;133;157m@[0m[38;2;140;131;156m@[0m[38;2;141;130;155m@[0m[38;2;136;120;149m@[0m[38;2;94;76;113m9[0m[38;2;83;66;99mS[0m[38;2;82;66;90mS[0m[38;2;95;78;94m#[0m[38;2;81;64;87mG[0m[38;2;80;63;98mS[0m[38;2;85;67;104m#[0m[38;2;79;63;93mS[0m[38;2;84;66;90mS[0m[38;2;83;62;81mG[0m[38;2;64;46;64mh[0m[38;2;56;38;57m5[0m[38;2;57;38;60m5[0m[38;2;55;39;60m5[0m[38;2;61;46;67mh[0m[38;2;69;54;73mM[0m[38;2;59;44;63m3[0m[38;2;51;37;58m5[0m[38;2;62;52;71mM[0m[38;2;87;71;88mS[0m[38;2;80;60;76mG[0m[38;2;53;36;55m5[0m[38;2;49;34;55m2[0m[38;2;48;35;56m2[0m[38;2;71;60;80mH[0m[38;2;95;78;96m#[0m[38;2;93;74;93m#[0m[38;2;96;77;96m#[0m[38;2;96;77;96m#[0m[38;2;83;63;76mG[0m[38;2;49;35;54m2[0m[38;2;72;60;82mH[0m[38;2;92;69;87mS[0m[38;2;65;51;67mh[0m[38;2;71;60;75mH[0m[38;2;50;46;61m3[0m[38;2;44;43;60m5[0m[38;2;44;43;59m5[0m[38;2;44;43;59m5[0m[38;2;44;43;59m5[0m[38;2;40;38;54m2[0m[38;2;39;37;55m2[0m[38;2;41;40;58m2[0m[38;2;45;44;62m5[0m[38;2;41;40;56m2[0m");
	$display("[38;2;149;130;149m@[0m[38;2;142;120;139m@[0m[38;2;142;117;136m@[0m[38;2;142;117;136m@[0m[38;2;143;117;138m@[0m[38;2;130;110;130m&[0m[38;2;133;113;131m&[0m[38;2;142;120;137m@[0m[38;2;140;119;137m@[0m[38;2;102;89;110m9[0m[38;2;112;89;105mB[0m[38;2;143;118;134m@[0m[38;2;142;117;136m@[0m[38;2;142;117;136m@[0m[38;2;149;128;143m@[0m[38;2;144;122;141m@[0m[38;2;142;117;135m@[0m[38;2;122;103;126m&[0m[38;2;76;60;88mG[0m[38;2;88;67;90mS[0m[38;2;99;81;102m9[0m[38;2;111;88;105mB[0m[38;2;145;124;138m@[0m[38;2;145;126;142m@[0m[38;2;140;116;134m@[0m[38;2;140;115;134m@[0m[38;2;140;115;134m@[0m[38;2;140;115;134m@[0m[38;2;139;116;135m@[0m[38;2;103;85;105m9[0m[38;2;123;98;117m&[0m[38;2;140;116;134m@[0m[38;2;141;120;137m@[0m[38;2;140;117;135m@[0m[38;2;139;114;133m@[0m[38;2;138;114;132m@[0m[38;2;135;112;131m&[0m[38;2;96;81;103m9[0m[38;2;70;52;77mH[0m[38;2;77;57;82mG[0m[38;2;76;56;83mH[0m[38;2;108;87;103m9[0m[38;2;116;96;113mB[0m[38;2;74;57;84mH[0m[38;2;84;64;93mS[0m[38;2;103;82;119mB[0m[38;2;101;82;121mB[0m[38;2;121;104;137m&[0m[38;2;157;146;166m@[0m[38;2;144;135;156m@[0m[38;2;116;99;116mB[0m[38;2;127;106;121m&[0m[38;2;105;84;107m9[0m[38;2;73;56;84mH[0m[38;2;88;69;101m#[0m[38;2;107;86;121mB[0m[38;2;137;122;148m@[0m[38;2;151;142;163m@[0m[38;2;150;143;163m@[0m[38;2;148;139;162m@[0m[38;2;120;106;125m&[0m[38;2;125;108;131m&[0m[38;2;106;88;124mB[0m[38;2;140;129;156m@[0m[38;2;146;139;162m@[0m[38;2;145;137;161m@[0m[38;2;145;137;161m@[0m[38;2;144;136;160m@[0m[38;2;139;131;155m@[0m[38;2;139;131;155m@[0m[38;2;141;133;157m@[0m[38;2;141;132;156m@[0m[38;2;134;120;148m@[0m[38;2;92;76;112m9[0m[38;2;90;68;107m#[0m[38;2;87;67;103m#[0m[38;2;80;63;91mS[0m[38;2;82;67;88mS[0m[38;2;79;63;84mG[0m[38;2;79;61;94mS[0m[38;2;82;65;102mS[0m[38;2;82;62;99mS[0m[38;2;80;61;90mG[0m[38;2;72;56;79mH[0m[38;2;62;47;66mh[0m[38;2;54;39;56m5[0m[38;2;52;37;57m5[0m[38;2;52;37;58m5[0m[38;2;53;38;59m5[0m[38;2;58;43;63m3[0m[38;2;56;41;62m3[0m[38;2;50;36;57m5[0m[38;2;55;40;61m3[0m[38;2;70;55;75mH[0m[38;2;67;51;68mM[0m[38;2;51;35;56m2[0m[38;2;48;33;54m2[0m[38;2;54;42;61m3[0m[38;2;88;71;92mS[0m[38;2;92;73;92m#[0m[38;2;94;74;94m#[0m[38;2;97;78;97m#[0m[38;2;92;71;88mS[0m[38;2;59;40;57m3[0m[38;2;55;45;64m3[0m[38;2;90;73;90mS[0m[38;2;73;55;68mM[0m[38;2;69;55;74mM[0m[38;2;60;49;64mh[0m[38;2;43;43;59m5[0m[38;2;42;41;57m2[0m[38;2;42;41;57m2[0m[38;2;42;41;57m2[0m[38;2;38;37;53mA[0m[38;2;38;37;54mA[0m[38;2;41;40;58m2[0m[38;2;45;44;61m5[0m[38;2;40;40;54m2[0m");
	$display("[38;2;149;129;148m@[0m[38;2;142;120;139m@[0m[38;2;142;117;136m@[0m[38;2;142;117;136m@[0m[38;2;142;118;136m@[0m[38;2;127;109;128m&[0m[38;2;122;100;119m&[0m[38;2;143;118;136m@[0m[38;2;142;119;137m@[0m[38;2;104;91;113mB[0m[38;2;102;80;98m9[0m[38;2;139;115;133m@[0m[38;2;141;117;136m@[0m[38;2;141;116;134m@[0m[38;2;148;128;142m@[0m[38;2;145;123;142m@[0m[38;2;141;116;135m@[0m[38;2;122;103;126m&[0m[38;2;76;59;87mG[0m[38;2;81;61;87mG[0m[38;2;89;68;90mS[0m[38;2;126;101;116m&[0m[38;2;147;127;140m@[0m[38;2;141;119;136m@[0m[38;2;139;116;134m@[0m[38;2;140;115;134m@[0m[38;2;140;115;134m@[0m[38;2;141;117;136m@[0m[38;2;113;95;117mB[0m[38;2;97;76;96m#[0m[38;2;139;113;131m@[0m[38;2;141;117;135m@[0m[38;2;140;120;137m@[0m[38;2;136;113;132m@[0m[38;2;136;111;129m&[0m[38;2;128;108;125m&[0m[38;2;94;77;98m#[0m[38;2;71;51;75mM[0m[38;2;84;65;90mS[0m[38;2;96;75;104m#[0m[38;2;103;79;103m9[0m[38;2;114;95;113mB[0m[38;2;73;58;84mH[0m[38;2;81;62;91mS[0m[38;2;103;81;115m9[0m[38;2;102;79;119m9[0m[38;2;123;104;134m&[0m[38;2;157;146;165m@[0m[38;2;147;138;155m@[0m[38;2;123;106;122m&[0m[38;2;127;105;120m&[0m[38;2;96;78;97m#[0m[38;2;76;57;84mG[0m[38;2;93;72;104m#[0m[38;2;111;92;124mB[0m[38;2;140;130;152m@[0m[38;2;151;142;162m@[0m[38;2;151;142;163m@[0m[38;2;151;143;164m@[0m[38;2;142;131;152m@[0m[38;2;119;104;122m&[0m[38;2;129;113;141m@[0m[38;2;106;91;124mB[0m[38;2;145;135;161m@[0m[38;2;146;138;162m@[0m[38;2;145;137;161m@[0m[38;2;145;137;161m@[0m[38;2;144;136;160m@[0m[38;2;141;133;157m@[0m[38;2;138;130;154m@[0m[38;2;141;133;157m@[0m[38;2;140;132;156m@[0m[38;2;133;123;149m@[0m[38;2;95;76;112m9[0m[38;2;88;67;105m#[0m[38;2;87;67;104m#[0m[38;2;81;65;99mS[0m[38;2;90;75;104m#[0m[38;2;93;78;99m#[0m[38;2;79;64;84mG[0m[38;2;73;57;82mH[0m[38;2;77;61;92mG[0m[38;2;102;87;120mB[0m[38;2;104;90;118mB[0m[38;2;80;66;92mS[0m[38;2;66;51;72mM[0m[38;2;56;41;62m3[0m[38;2;53;38;59m5[0m[38;2;52;37;58m5[0m[38;2;51;36;57m5[0m[38;2;52;36;58m5[0m[38;2;51;36;57m5[0m[38;2;50;35;56m2[0m[38;2;49;33;54m2[0m[38;2;52;37;58m5[0m[38;2;53;34;56m5[0m[38;2;52;33;54m2[0m[38;2;49;33;53m2[0m[38;2;72;57;79mH[0m[38;2;86;67;85mS[0m[38;2;87;69;87mS[0m[38;2;96;77;96m#[0m[38;2;95;74;92m#[0m[38;2;74;53;67mM[0m[38;2;45;34;51mA[0m[38;2;78;63;85mG[0m[38;2;87;66;81mS[0m[38;2;60;45;61m3[0m[38;2;74;57;75mH[0m[38;2;46;43;57m5[0m[38;2;42;41;57m2[0m[38;2;42;41;57m2[0m[38;2;40;39;55m2[0m[38;2;36;35;51mA[0m[38;2;37;36;52mA[0m[38;2;41;40;56m2[0m[38;2;43;41;58m2[0m[38;2;38;38;52mA[0m");
	$display("[38;2;149;128;145m@[0m[38;2;141;119;136m@[0m[38;2;142;116;135m@[0m[38;2;140;116;134m@[0m[38;2;134;113;130m&[0m[38;2;126;110;128m&[0m[38;2;110;90;110mB[0m[38;2;141;116;132m@[0m[38;2;142;117;138m@[0m[38;2;108;94;117mB[0m[38;2;92;72;94m#[0m[38;2;137;112;130m@[0m[38;2;141;116;135m@[0m[38;2;140;115;134m@[0m[38;2;148;127;141m@[0m[38;2;144;123;143m@[0m[38;2;141;116;137m@[0m[38;2;124;104;128m&[0m[38;2;76;60;86mG[0m[38;2;72;53;80mH[0m[38;2;83;62;83mG[0m[38;2;135;110;125m&[0m[38;2;146;124;137m@[0m[38;2;140;115;134m@[0m[38;2;140;115;134m@[0m[38;2;140;115;134m@[0m[38;2;141;116;135m@[0m[38;2;124;106;127m&[0m[38;2;85;67;88mS[0m[38;2;126;100;116m&[0m[38;2;139;114;129m@[0m[38;2;137;114;129m@[0m[38;2;130;108;124m&[0m[38;2;131;108;124m&[0m[38;2;128;105;123m&[0m[38;2;92;75;97m#[0m[38;2;70;52;78mH[0m[38;2;87;68;92mS[0m[38;2;98;79;110m9[0m[38;2;95;76;97m#[0m[38;2;103;87;105m9[0m[38;2;75;56;81mH[0m[38;2;81;61;88mG[0m[38;2;102;80;115m9[0m[38;2;103;81;118m9[0m[38;2;126;108;139m&[0m[38;2;158;148;166m@[0m[38;2;146;137;152m@[0m[38;2;127;108;124m&[0m[38;2;121;101;117m&[0m[38;2;86;71;92mS[0m[38;2;78;62;88mG[0m[38;2;95;76;110m9[0m[38;2;119;99;129m&[0m[38;2;147;135;156m@[0m[38;2;151;143;161m@[0m[38;2;153;144;162m@[0m[38;2;151;142;161m@[0m[38;2;153;143;164m@[0m[38;2;128;116;137m@[0m[38;2;132;117;139m@[0m[38;2;122;106;138m&[0m[38;2;114;99;130m&[0m[38;2;149;138;163m@[0m[38;2;146;138;162m@[0m[38;2;145;137;161m@[0m[38;2;145;137;161m@[0m[38;2;145;137;161m@[0m[38;2;143;135;159m@[0m[38;2;138;130;154m@[0m[38;2;140;131;156m@[0m[38;2;140;132;156m@[0m[38;2;136;125;150m@[0m[38;2;97;78;112m9[0m[38;2;86;68;105m#[0m[38;2;82;66;100mS[0m[38;2;100;88;116mB[0m[38;2;118;107;132m&[0m[38;2;106;99;120mB[0m[38;2;74;64;82mG[0m[38;2;51;40;57m5[0m[38;2;54;42;61m3[0m[38;2;58;46;67mh[0m[38;2;68;59;79mH[0m[38;2;81;68;89mS[0m[38;2;76;59;79mH[0m[38;2;63;48;67mh[0m[38;2;54;40;59m5[0m[38;2;48;34;54m2[0m[38;2;48;35;55m2[0m[38;2;50;36;56m2[0m[38;2;51;36;57m5[0m[38;2;51;34;55m2[0m[38;2;51;33;54m2[0m[38;2;51;32;54m2[0m[38;2;51;32;54m2[0m[38;2;51;33;54m2[0m[38;2;47;31;52mA[0m[38;2;54;43;62m3[0m[38;2;86;67;85mS[0m[38;2;74;58;75mH[0m[38;2;91;75;94m#[0m[38;2;95;75;92m#[0m[38;2;84;63;79mG[0m[38;2;47;32;49mA[0m[38;2;63;49;71mh[0m[38;2;92;70;86mS[0m[38;2;63;44;58m3[0m[38;2;69;54;74mM[0m[38;2;58;45;61m3[0m[38;2;43;42;55m2[0m[38;2;42;40;56m2[0m[38;2;39;36;53mA[0m[38;2;37;34;51mA[0m[38;2;38;35;52mA[0m[38;2;41;38;55m2[0m[38;2;42;39;56m2[0m[38;2;37;34;50mA[0m");
	$display("[38;2;148;128;144m@[0m[38;2;140;118;135m@[0m[38;2;141;115;134m@[0m[38;2;138;114;132m@[0m[38;2;129;107;124m&[0m[38;2;132;112;132m&[0m[38;2;100;83;103m9[0m[38;2;134;109;124m&[0m[38;2;142;118;135m@[0m[38;2;114;99;118mB[0m[38;2;86;67;91mS[0m[38;2;132;108;123m&[0m[38;2;141;116;135m@[0m[38;2;140;115;133m@[0m[38;2;145;124;137m@[0m[38;2;146;126;143m@[0m[38;2;142;116;135m@[0m[38;2;125;105;125m&[0m[38;2;76;61;85mG[0m[38;2;70;54;79mH[0m[38;2;88;66;85mS[0m[38;2;141;114;129m@[0m[38;2;141;120;135m@[0m[38;2;140;115;134m@[0m[38;2;139;115;134m@[0m[38;2;138;114;132m@[0m[38;2;132;110;128m&[0m[38;2;85;68;93mS[0m[38;2;102;78;97m9[0m[38;2;133;108;122m&[0m[38;2;135;111;125m&[0m[38;2;134;110;125m&[0m[38;2;135;112;127m&[0m[38;2;130;109;125m&[0m[38;2;90;75;97m#[0m[38;2;71;53;77mH[0m[38;2;90;70;97m#[0m[38;2;101;82;114m9[0m[38;2;90;72;98m#[0m[38;2;91;73;93m#[0m[38;2;72;55;76mH[0m[38;2;86;64;89mS[0m[38;2;104;81;114m9[0m[38;2;108;86;120mB[0m[38;2;136;120;145m@[0m[38;2;159;150;168m@[0m[38;2;146;135;153m@[0m[38;2;128;110;126m&[0m[38;2;109;88;107mB[0m[38;2;82;65;87mS[0m[38;2;86;68;100m#[0m[38;2;104;82;116m9[0m[38;2;130;112;140m@[0m[38;2;152;141;161m@[0m[38;2;151;143;161m@[0m[38;2;153;144;164m@[0m[38;2;153;144;164m@[0m[38;2;153;144;164m@[0m[38;2;145;133;155m@[0m[38;2;122;107;130m&[0m[38;2;148;133;159m@[0m[38;2;107;91;125mB[0m[38;2;131;118;148m@[0m[38;2;148;138;163m@[0m[38;2;146;137;161m@[0m[38;2;145;137;161m@[0m[38;2;145;137;161m@[0m[38;2;144;136;160m@[0m[38;2;142;135;158m@[0m[38;2;139;133;156m@[0m[38;2;138;129;153m@[0m[38;2;140;132;156m@[0m[38;2;138;130;154m@[0m[38;2;103;87;118mB[0m[38;2;87;69;105m#[0m[38;2;116;102;133m&[0m[38;2;128;116;139m@[0m[38;2;83;72;87mS[0m[38;2;48;37;49m2[0m[38;2;40;31;42mX[0m[38;2;38;32;42mX[0m[38;2;40;33;45mX[0m[38;2;49;41;53m5[0m[38;2;50;39;55m5[0m[38;2;58;45;62m3[0m[38;2;58;42;57m3[0m[38;2;46;33;43mA[0m[38;2;39;28;37ms[0m[38;2;33;25;34mr[0m[38;2;32;25;35mr[0m[38;2;34;28;40ms[0m[38;2;43;34;49mA[0m[38;2;51;36;58m5[0m[38;2;56;38;61m5[0m[38;2;54;35;57m5[0m[38;2;51;32;54m2[0m[38;2;50;32;54m2[0m[38;2;46;31;52mA[0m[38;2;45;34;53m2[0m[38;2;77;61;79mG[0m[38;2;70;52;69mM[0m[38;2;84;70;92mS[0m[38;2;93;76;93m#[0m[38;2;91;69;84mS[0m[38;2;54;37;50m2[0m[38;2;48;38;57m5[0m[38;2;85;70;86mS[0m[38;2;76;54;66mM[0m[38;2;56;43;62m3[0m[38;2;71;55;71mM[0m[38;2;41;38;55m2[0m[38;2;41;38;55m2[0m[38;2;36;33;50mA[0m[38;2;35;32;49mX[0m[38;2;36;33;50mA[0m[38;2;40;37;54m2[0m[38;2;40;38;54m2[0m[38;2;35;34;49mX[0m");
	$display("[38;2;148;127;144m@[0m[38;2;141;119;136m@[0m[38;2;141;115;134m@[0m[38;2;136;113;133m@[0m[38;2;126;102;121m&[0m[38;2;136;113;131m@[0m[38;2;96;78;101m#[0m[38;2;119;95;113mB[0m[38;2;143;118;132m@[0m[38;2;122;104;124m&[0m[38;2;81;65;89mS[0m[38;2;126;101;115m&[0m[38;2;141;117;134m@[0m[38;2;140;115;134m@[0m[38;2;142;120;135m@[0m[38;2;145;127;142m@[0m[38;2;140;117;135m@[0m[38;2;127;107;126m&[0m[38;2;78;63;87mG[0m[38;2;71;52;78mH[0m[38;2;90;67;87mS[0m[38;2;141;115;129m@[0m[38;2;137;114;130m@[0m[38;2;134;109;127m&[0m[38;2;132;107;124m&[0m[38;2;128;108;124m&[0m[38;2;89;75;95m#[0m[38;2;90;67;87mS[0m[38;2;137;110;124m&[0m[38;2;141;115;129m@[0m[38;2;141;116;130m@[0m[38;2;140;116;132m@[0m[38;2;126;107;125m&[0m[38;2;86;68;91mS[0m[38;2;71;54;78mH[0m[38;2;94;75;102m#[0m[38;2;101;80;114m9[0m[38;2;79;64;90mG[0m[38;2;76;61;80mG[0m[38;2;73;54;76mH[0m[38;2;90;69;98m#[0m[38;2;102;80;115m9[0m[38;2;106;86;119mB[0m[38;2;134;117;144m@[0m[38;2;150;138;160m@[0m[38;2;140;127;146m@[0m[38;2;117;97;116mB[0m[38;2;93;74;94m#[0m[38;2;85;65;96mS[0m[38;2;98;76;112m9[0m[38;2;116;97;129m&[0m[38;2;144;131;153m@[0m[38;2;155;146;163m@[0m[38;2;152;143;162m@[0m[38;2;153;144;167m@[0m[38;2;153;144;165m@[0m[38;2;153;145;165m@[0m[38;2;151;141;163m@[0m[38;2;125;112;134m&[0m[38;2;144;130;154m@[0m[38;2;137;123;150m@[0m[38;2;109;95;126mB[0m[38;2;145;136;161m@[0m[38;2;146;137;161m@[0m[38;2;146;136;161m@[0m[38;2;145;137;161m@[0m[38;2;145;137;161m@[0m[38;2;144;136;160m@[0m[38;2;142;134;158m@[0m[38;2;142;134;158m@[0m[38;2;138;130;154m@[0m[38;2;137;129;153m@[0m[38;2;139;131;155m@[0m[38;2;129;118;144m@[0m[38;2;117;105;131m&[0m[38;2;118;108;127m&[0m[38;2;84;71;85mS[0m[38;2;58;45;55m3[0m[38;2;57;46;60m3[0m[38;2;61;57;79mM[0m[38;2;65;63;94mG[0m[38;2;67;65;99mG[0m[38;2;69;67;101mS[0m[38;2;68;67;100mS[0m[38;2;64;63;94mG[0m[38;2;59;56;82mM[0m[38;2;57;52;72mh[0m[38;2;54;48;69mh[0m[38;2;49;43;60m5[0m[38;2;39;35;44mX[0m[38;2;30;27;32mr[0m[38;2;28;22;27mi[0m[38;2;34;29;43ms[0m[38;2;52;43;64m3[0m[38;2;55;42;65m3[0m[38;2;60;42;68mh[0m[38;2;66;48;74mM[0m[38;2;57;42;63m3[0m[38;2;44;30;49mA[0m[38;2;66;50;70mM[0m[38;2;69;51;66mM[0m[38;2;74;61;80mH[0m[38;2;92;75;93m#[0m[38;2;93;70;88mS[0m[38;2;64;44;58m3[0m[38;2;42;30;50mA[0m[38;2;75;61;79mH[0m[38;2;85;63;76mG[0m[38;2;51;35;52m2[0m[38;2;72;57;74mH[0m[38;2;50;41;56m5[0m[38;2;40;38;54m2[0m[38;2;35;32;48mX[0m[38;2;35;32;49mX[0m[38;2;36;33;50mA[0m[38;2;37;34;52mA[0m[38;2;37;35;52mA[0m[38;2;34;33;48mX[0m");
	$display("[38;2;147;126;142m@[0m[38;2;140;118;136m@[0m[38;2;140;115;134m@[0m[38;2;135;113;133m@[0m[38;2;117;96;116mB[0m[38;2;136;113;129m&[0m[38;2;96;81;106m9[0m[38;2;98;76;96m#[0m[38;2;140;115;128m@[0m[38;2;129;110;129m&[0m[38;2;81;67;92mS[0m[38;2;117;90;107mB[0m[38;2;141;116;133m@[0m[38;2;140;115;134m@[0m[38;2;141;116;135m@[0m[38;2;147;125;143m@[0m[38;2;140;117;135m@[0m[38;2;130;110;129m&[0m[38;2;80;65;90mS[0m[38;2;70;52;78mH[0m[38;2;88;65;85mS[0m[38;2;131;107;121m&[0m[38;2;132;108;122m&[0m[38;2;135;111;124m&[0m[38;2;137;114;128m@[0m[38;2;100;86;107m9[0m[38;2;78;61;80mG[0m[38;2;129;103;116m&[0m[38;2;141;116;130m@[0m[38;2;139;115;129m@[0m[38;2;140;116;129m@[0m[38;2;118;99;116mB[0m[38;2;77;62;83mG[0m[38;2;76;57;82mH[0m[38;2;99;78;106m9[0m[38;2;97;77;111m9[0m[38;2;76;57;86mG[0m[38;2;70;53;76mH[0m[38;2;77;59;83mG[0m[38;2;93;72;101m#[0m[38;2;103;84;117mB[0m[38;2;109;93;125mB[0m[38;2;106;91;123mB[0m[38;2;105;89;117mB[0m[38;2;110;91;113mB[0m[38;2;96;76;99m#[0m[38;2;85;65;95mS[0m[38;2;95;73;110m9[0m[38;2;113;93;126mB[0m[38;2;137;123;148m@[0m[38;2;155;145;164m@[0m[38;2;154;146;164m@[0m[38;2;153;144;163m@[0m[38;2;155;146;166m@[0m[38;2;153;143;167m@[0m[38;2;154;145;165m@[0m[38;2;152;141;162m@[0m[38;2;130;119;138m@[0m[38;2;140;129;148m@[0m[38;2;151;138;164m@[0m[38;2;115;100;129m&[0m[38;2;137;124;153m@[0m[38;2;148;138;163m@[0m[38;2;146;136;161m@[0m[38;2;146;136;161m@[0m[38;2;145;137;160m@[0m[38;2;144;136;159m@[0m[38;2;144;136;160m@[0m[38;2;142;134;158m@[0m[38;2;141;133;157m@[0m[38;2;141;133;157m@[0m[38;2;136;128;152m@[0m[38;2;137;129;153m@[0m[38;2;138;130;154m@[0m[38;2;128;120;142m@[0m[38;2;107;96;114mB[0m[38;2;72;57;71mH[0m[38;2;64;57;77mM[0m[38;2;64;63;95mG[0m[38;2;69;70;107mS[0m[38;2;72;72;108mS[0m[38;2;73;73;108m#[0m[38;2;59;59;92mH[0m[38;2;53;55;84mM[0m[38;2;53;54;84mM[0m[38;2;54;55;87mM[0m[38;2;53;55;84mM[0m[38;2;56;57;88mH[0m[38;2;65;64;96mG[0m[38;2;64;60;91mH[0m[38;2;59;55;80mM[0m[38;2;48;43;61m5[0m[38;2;33;29;35mr[0m[38;2;26;21;26m;[0m[38;2;32;26;38mr[0m[38;2;52;44;65m3[0m[38;2;68;54;82mH[0m[38;2;61;46;67mh[0m[38;2;44;30;47mA[0m[38;2;56;40;61m3[0m[38;2;67;50;67mM[0m[38;2;65;52;69mM[0m[38;2;92;73;91m#[0m[38;2;93;69;88mS[0m[38;2;73;51;65mM[0m[38;2;41;26;47mX[0m[38;2;61;50;70mh[0m[38;2;87;68;83mS[0m[38;2;55;37;51m5[0m[38;2;61;50;69mh[0m[38;2;63;48;60mh[0m[38;2;34;32;44mX[0m[38;2;33;31;45mX[0m[38;2;30;28;45ms[0m[38;2;34;32;48mX[0m[38;2;35;33;50mX[0m[38;2;35;33;50mX[0m[38;2;33;31;46mX[0m");
	$display("[38;2;147;127;141m@[0m[38;2;140;118;137m@[0m[38;2;141;115;134m@[0m[38;2;135;113;131m@[0m[38;2;110;91;111mB[0m[38;2;135;112;127m&[0m[38;2;100;88;111m9[0m[38;2;80;62;83mG[0m[38;2;129;103;115m&[0m[38;2;135;116;131m@[0m[38;2;87;73;97m#[0m[38;2;106;80;99m9[0m[38;2;141;115;130m@[0m[38;2;140;115;132m@[0m[38;2;139;115;132m@[0m[38;2;147;122;138m@[0m[38;2;142;117;133m@[0m[38;2;133;113;129m&[0m[38;2;83;69;93mS[0m[38;2;69;50;73mM[0m[38;2;86;64;82mG[0m[38;2;136;110;125m&[0m[38;2;142;116;129m@[0m[38;2;140;117;133m@[0m[38;2;107;89;112mB[0m[38;2;75;57;79mH[0m[38;2;121;95;110mB[0m[38;2;140;115;129m@[0m[38;2;140;115;129m@[0m[38;2;135;114;128m&[0m[38;2;105;88;108m9[0m[38;2;72;57;79mH[0m[38;2;84;62;89mS[0m[38;2;102;81;113m9[0m[38;2;90;72;104m#[0m[38;2;72;55;81mH[0m[38;2;75;58;79mH[0m[38;2;92;71;97m#[0m[38;2;103;81;115m9[0m[38;2;115;97;126m&[0m[38;2;146;131;152m@[0m[38;2;153;139;159m@[0m[38;2;123;109;130m&[0m[38;2;91;75;96m#[0m[38;2;83;65;90mS[0m[38;2;99;78;108m9[0m[38;2;117;97;128m&[0m[38;2;137;122;148m@[0m[38;2;156;146;166m@[0m[38;2;157;149;167m@[0m[38;2;153;144;163m@[0m[38;2;154;145;164m@[0m[38;2;155;146;166m@[0m[38;2;156;147;167m@[0m[38;2;154;145;165m@[0m[38;2;145;136;156m@[0m[38;2;133;121;142m@[0m[38;2;146;132;152m@[0m[38;2;153;141;163m@[0m[38;2;128;115;141m@[0m[38;2;135;122;149m@[0m[38;2;150;138;164m@[0m[38;2;146;136;161m@[0m[38;2;146;136;161m@[0m[38;2;146;136;161m@[0m[38;2;145;137;158m@[0m[38;2;144;135;156m@[0m[38;2;143;135;157m@[0m[38;2;142;134;157m@[0m[38;2;141;133;157m@[0m[38;2;141;133;157m@[0m[38;2;139;131;155m@[0m[38;2;135;127;151m@[0m[38;2;137;129;153m@[0m[38;2;132;123;146m@[0m[38;2;104;94;111mB[0m[38;2;94;85;108m9[0m[38;2;72;72;108mS[0m[38;2;84;84;122m9[0m[38;2;105;102;138m&[0m[38;2;115;111;146m&[0m[38;2;64;63;91mG[0m[38;2;44;45;74m3[0m[38;2;47;48;78mh[0m[38;2;42;44;72m3[0m[38;2;38;40;66m5[0m[38;2;36;37;63m2[0m[38;2;31;33;58mA[0m[38;2;56;61;92mH[0m[38;2;93;92;126mB[0m[38;2;84;79;112m#[0m[38;2;67;64;100mG[0m[38;2;60;58;85mH[0m[38;2;41;38;51mA[0m[38;2;28;21;28mi[0m[38;2;28;22;30mi[0m[38;2;46;36;59m2[0m[38;2;57;44;65m3[0m[38;2;45;29;48mA[0m[38;2;48;35;55m2[0m[38;2;64;47;62mh[0m[38;2;57;44;63m3[0m[38;2;89;71;90mS[0m[38;2;92;70;88mS[0m[38;2;80;58;72mH[0m[38;2;43;27;46mX[0m[38;2;50;39;60m5[0m[38;2;86;67;83mS[0m[38;2;64;44;57m3[0m[38;2;48;38;57m5[0m[38;2;73;57;71mH[0m[38;2;36;32;44mX[0m[38;2;34;34;49mX[0m[38;2;33;31;47mX[0m[38;2;32;30;47mX[0m[38;2;31;30;46ms[0m[38;2;31;30;46ms[0m[38;2;29;28;42ms[0m");
	$display("[38;2;146;126;140m@[0m[38;2;140;118;137m@[0m[38;2;141;115;134m@[0m[38;2;135;113;131m@[0m[38;2;104;86;106m9[0m[38;2;131;108;122m&[0m[38;2;107;94;116mB[0m[38;2;72;56;80mH[0m[38;2;110;84;97m9[0m[38;2;139;116;129m@[0m[38;2;98;83;104m9[0m[38;2;94;73;90m#[0m[38;2;139;113;126m&[0m[38;2;139;115;129m@[0m[38;2;139;115;129m@[0m[38;2;144;120;133m@[0m[38;2;142;119;132m@[0m[38;2;137;114;129m@[0m[38;2;88;75;97m#[0m[38;2;68;52;73mM[0m[38;2;83;61;82mG[0m[38;2;134;107;123m&[0m[38;2;141;115;130m@[0m[38;2;108;91;112mB[0m[38;2;75;57;81mH[0m[38;2;116;91;106mB[0m[38;2;141;114;128m@[0m[38;2;139;115;129m@[0m[38;2;127;106;122m&[0m[38;2;90;73;94m#[0m[38;2;73;55;79mH[0m[38;2;90;70;97m#[0m[38;2;97;75;106m9[0m[38;2;80;60;91mG[0m[38;2;69;52;74mM[0m[38;2;79;61;83mG[0m[38;2;83;68;91mS[0m[38;2;76;64;86mG[0m[38;2;69;58;79mH[0m[38;2;85;74;89mS[0m[38;2;99;85;101m9[0m[38;2;86;73;91mS[0m[38;2;71;55;71mM[0m[38;2;73;55;71mH[0m[38;2;91;73;93m#[0m[38;2;120;108;125m&[0m[38;2;142;133;150m@[0m[38;2;146;139;155m@[0m[38;2;145;137;154m@[0m[38;2;150;141;160m@[0m[38;2;155;146;165m@[0m[38;2;155;146;165m@[0m[38;2;154;145;164m@[0m[38;2;148;139;158m@[0m[38;2;138;129;148m@[0m[38;2;138;129;147m@[0m[38;2;149;139;159m@[0m[38;2;150;139;161m@[0m[38;2;138;127;152m@[0m[38;2;142;132;157m@[0m[38;2;150;141;166m@[0m[38;2;147;138;163m@[0m[38;2;146;136;161m@[0m[38;2;146;136;161m@[0m[38;2;146;136;161m@[0m[38;2;145;136;158m@[0m[38;2;144;135;156m@[0m[38;2;142;134;155m@[0m[38;2;141;133;155m@[0m[38;2;141;133;157m@[0m[38;2;141;133;157m@[0m[38;2;140;132;156m@[0m[38;2;137;129;153m@[0m[38;2;136;128;152m@[0m[38;2;128;120;143m@[0m[38;2;128;119;140m@[0m[38;2;127;120;146m@[0m[38;2;114;111;146m&[0m[38;2;132;128;163m@[0m[38;2;137;131;167m@[0m[38;2;127;122;153m@[0m[38;2;82;78;102m#[0m[38;2;76;75;99mS[0m[38;2;45;44;66m5[0m[38;2;31;32;53mX[0m[38;2;47;49;71m3[0m[38;2;40;42;65m5[0m[38;2;43;44;70m3[0m[38;2;39;42;68m5[0m[38;2;63;67;98mG[0m[38;2;116;115;150m@[0m[38;2;103;96;129mB[0m[38;2;70;68;101mS[0m[38;2;64;60;94mG[0m[38;2;51;45;66m3[0m[38;2;32;26;31mr[0m[38;2;29;23;29mi[0m[38;2;34;28;39ms[0m[38;2;42;31;48mA[0m[38;2;44;31;49mA[0m[38;2;55;40;55m5[0m[38;2;51;40;57m5[0m[38;2;88;70;88mS[0m[38;2;93;69;88mS[0m[38;2;84;63;76mG[0m[38;2;47;30;45mA[0m[38;2;44;32;52mA[0m[38;2;79;63;80mG[0m[38;2;73;52;65mM[0m[38;2;42;30;46mX[0m[38;2;74;59;74mH[0m[38;2;53;39;52m5[0m[38;2;35;33;50mX[0m[38;2;37;34;52mA[0m[38;2;34;31;48mX[0m[38;2;34;32;48mX[0m[38;2;33;31;46mX[0m[38;2;29;28;40mr[0m");
	$display("[38;2;145;125;139m@[0m[38;2;140;118;137m@[0m[38;2;140;115;134m@[0m[38;2;135;113;131m@[0m[38;2;99;81;104m9[0m[38;2;126;100;115m&[0m[38;2;114;99;119mB[0m[38;2;70;58;82mH[0m[38;2;87;65;83mS[0m[38;2;134;109;122m&[0m[38;2;111;94;113mB[0m[38;2;86;68;86mS[0m[38;2;135;109;122m&[0m[38;2;140;116;130m@[0m[38;2;139;115;129m@[0m[38;2;140;117;131m@[0m[38;2;143;122;134m@[0m[38;2;138;116;130m@[0m[38;2;99;85;105m9[0m[38;2;66;53;75mM[0m[38;2;78;56;78mH[0m[38;2;128;102;117m&[0m[38;2;107;91;111mB[0m[38;2;74;58;80mH[0m[38;2;116;89;106mB[0m[38;2;142;114;129m@[0m[38;2;136;111;126m&[0m[38;2;109;90;108mB[0m[38;2;78;61;84mG[0m[38;2;80;61;85mG[0m[38;2;92;72;98m#[0m[38;2;85;63;93mS[0m[38;2;78;57;79mH[0m[38;2;84;63;81mG[0m[38;2;94;70;88mS[0m[38;2;99;74;91m#[0m[38;2;75;58;72mH[0m[38;2;61;49;59m3[0m[38;2;69;57;68mM[0m[38;2;68;56;68mM[0m[38;2;62;50;64mh[0m[38;2;63;51;65mh[0m[38;2;68;54;68mM[0m[38;2;75;57;71mH[0m[38;2;81;61;73mH[0m[38;2;86;65;77mG[0m[38;2;99;83;94m9[0m[38;2;114;102;115mB[0m[38;2;134;122;138m@[0m[38;2;146;136;155m@[0m[38;2;151;142;162m@[0m[38;2;153;144;163m@[0m[38;2;149;140;159m@[0m[38;2;147;138;157m@[0m[38;2;148;139;158m@[0m[38;2;148;139;158m@[0m[38;2;147;138;157m@[0m[38;2;147;138;158m@[0m[38;2;149;141;163m@[0m[38;2;149;141;164m@[0m[38;2;148;140;164m@[0m[38;2;147;138;163m@[0m[38;2;146;136;161m@[0m[38;2;146;136;161m@[0m[38;2;146;136;161m@[0m[38;2;145;136;158m@[0m[38;2;144;135;156m@[0m[38;2;143;134;155m@[0m[38;2;142;134;156m@[0m[38;2;140;132;156m@[0m[38;2;140;132;156m@[0m[38;2;139;131;155m@[0m[38;2;138;130;154m@[0m[38;2;137;130;154m@[0m[38;2;136;128;152m@[0m[38;2;136;128;151m@[0m[38;2;135;127;153m@[0m[38;2;137;130;164m@[0m[38;2;135;129;165m@[0m[38;2;136;130;165m@[0m[38;2;135;130;159m@[0m[38;2;105;104;131m&[0m[38;2;81;80;107m#[0m[38;2;56;57;86mH[0m[38;2;45;47;75m3[0m[38;2;54;58;92mH[0m[38;2;64;69;105mS[0m[38;2;47;51;76mh[0m[38;2;42;45;72m3[0m[38;2;34;39;67m2[0m[38;2;88;92;128mB[0m[38;2;125;119;157m@[0m[38;2;106;102;134m&[0m[38;2;67;65;98mG[0m[38;2;61;59;93mH[0m[38;2;47;41;53m2[0m[38;2;42;32;43mX[0m[38;2;54;42;61m3[0m[38;2;44;31;49mA[0m[38;2;42;29;45mX[0m[38;2;45;30;49mA[0m[38;2;48;37;55m2[0m[38;2;85;68;86mS[0m[38;2;93;68;88mS[0m[38;2;88;64;79mG[0m[38;2;52;33;46m2[0m[38;2;40;26;47mX[0m[38;2;71;57;75mH[0m[38;2;81;58;71mH[0m[38;2;44;28;46mX[0m[38;2;65;53;71mM[0m[38;2;67;49;61mh[0m[38;2;32;31;45mX[0m[38;2;37;35;49mA[0m[38;2;35;32;48mX[0m[38;2;35;32;49mX[0m[38;2;35;32;48mX[0m[38;2;31;29;43ms[0m");
	$display("[38;2;143;122;137m@[0m[38;2;140;117;137m@[0m[38;2;139;114;133m@[0m[38;2;135;113;131m@[0m[38;2;93;79;102m#[0m[38;2;116;92;107mB[0m[38;2;121;101;121m&[0m[38;2;73;60;85mG[0m[38;2;74;54;75mH[0m[38;2;117;92;105mB[0m[38;2;124;105;123m&[0m[38;2;84;67;87mS[0m[38;2;129;103;117m&[0m[38;2;142;115;130m@[0m[38;2;139;115;129m@[0m[38;2;139;116;129m@[0m[38;2;143;120;134m@[0m[38;2;139;116;129m@[0m[38;2;110;95;114mB[0m[38;2;69;54;77mH[0m[38;2;74;53;75mH[0m[38;2;88;69;89mS[0m[38;2;75;56;76mH[0m[38;2;115;89;105mB[0m[38;2;137;111;125m&[0m[38;2;114;94;112mB[0m[38;2;86;69;90mS[0m[38;2;76;58;83mG[0m[38;2;81;62;88mG[0m[38;2;76;59;80mH[0m[38;2;63;48;67mh[0m[38;2;59;46;62m3[0m[38;2;62;48;61mh[0m[38;2;71;56;69mM[0m[38;2;83;66;84mG[0m[38;2;87;71;94mS[0m[38;2;84;75;100m#[0m[38;2;82;75;104m#[0m[38;2;82;78;112m#[0m[38;2;82;81;115m9[0m[38;2;84;82;118m9[0m[38;2;83;81;118m9[0m[38;2;80;79;111m#[0m[38;2;78;75;106m#[0m[38;2;77;72;101mS[0m[38;2;80;72;99mS[0m[38;2;94;81;100m#[0m[38;2;101;86;99m9[0m[38;2;106;92;107mB[0m[38;2;122;109;128m&[0m[38;2;140;128;148m@[0m[38;2;150;140;160m@[0m[38;2;155;146;165m@[0m[38;2;155;146;165m@[0m[38;2;152;143;162m@[0m[38;2;151;142;161m@[0m[38;2;150;141;160m@[0m[38;2;150;141;160m@[0m[38;2;149;141;162m@[0m[38;2;149;141;162m@[0m[38;2;147;139;163m@[0m[38;2;146;138;162m@[0m[38;2;147;137;162m@[0m[38;2;146;136;161m@[0m[38;2;146;136;161m@[0m[38;2;145;137;159m@[0m[38;2;145;135;157m@[0m[38;2;144;134;155m@[0m[38;2;141;133;155m@[0m[38;2;140;131;156m@[0m[38;2;139;130;154m@[0m[38;2;139;129;154m@[0m[38;2;138;129;154m@[0m[38;2;138;130;154m@[0m[38;2;137;128;152m@[0m[38;2;134;126;151m@[0m[38;2;134;126;151m@[0m[38;2;134;127;157m@[0m[38;2;134;129;162m@[0m[38;2;134;128;164m@[0m[38;2;121;116;148m@[0m[38;2;48;47;70m3[0m[38;2;37;40;66m5[0m[38;2;58;67;105mG[0m[38;2;65;72;114mS[0m[38;2;56;63;106mG[0m[38;2;73;79;132m9[0m[38;2;63;70;111mS[0m[38;2;62;67;111mS[0m[38;2;61;66;104mG[0m[38;2;71;77;110m#[0m[38;2;122;116;155m@[0m[38;2;122;115;152m@[0m[38;2;88;83;115m9[0m[38;2;58;60;90mH[0m[38;2;52;45;63m3[0m[38;2;58;45;67mh[0m[38;2;68;52;79mH[0m[38;2;47;33;49mA[0m[38;2;43;29;46mX[0m[38;2;42;27;47mX[0m[38;2;46;34;54m2[0m[38;2;83;66;85mS[0m[38;2;93;68;88mS[0m[38;2;90;64;81mS[0m[38;2;55;36;49m2[0m[38;2;39;25;43ms[0m[38;2;63;50;67mh[0m[38;2;84;63;73mG[0m[38;2;46;30;44mA[0m[38;2;57;45;64m3[0m[38;2;78;58;70mH[0m[38;2;38;32;45mX[0m[38;2;33;32;48mX[0m[38;2;36;34;50mA[0m[38;2;35;32;49mX[0m[38;2;35;32;49mX[0m[38;2;31;29;44ms[0m");
	$display("[38;2;141;120;132m@[0m[38;2;140;118;134m@[0m[38;2;139;115;130m@[0m[38;2;136;115;130m@[0m[38;2;93;81;102m9[0m[38;2;104;79;96m9[0m[38;2;123;103;122m&[0m[38;2;76;63;87mG[0m[38;2;71;52;76mH[0m[38;2;94;70;87mS[0m[38;2;130;109;123m&[0m[38;2;90;74;94m#[0m[38;2;121;96;107mB[0m[38;2;141;114;129m@[0m[38;2;136;112;126m&[0m[38;2;135;111;125m&[0m[38;2;141;117;131m@[0m[38;2;141;117;129m@[0m[38;2;121;105;120m&[0m[38;2;74;57;81mH[0m[38;2;70;50;74mM[0m[38;2;71;52;73mM[0m[38;2;99;78;92m#[0m[38;2;108;88;104m9[0m[38;2;84;64;86mS[0m[38;2;71;53;75mH[0m[38;2;70;53;74mM[0m[38;2;66;51;70mM[0m[38;2;57;44;60m3[0m[38;2;51;39;52m2[0m[38;2;50;38;52m2[0m[38;2;57;46;62m3[0m[38;2;71;64;85mG[0m[38;2;81;76;105m#[0m[38;2;86;82;119m9[0m[38;2;85;84;124m9[0m[38;2;80;80;119m9[0m[38;2;77;78;116m#[0m[38;2;77;77;115m#[0m[38;2;78;78;117m#[0m[38;2;79;80;118m9[0m[38;2;92;92;130mB[0m[38;2;104;104;142m&[0m[38;2;103;105;143m&[0m[38;2;102;102;141m&[0m[38;2;98;99;138m&[0m[38;2;97;98;134mB[0m[38;2;122;117;146m@[0m[38;2;150;138;160m@[0m[38;2;147;134;153m@[0m[38;2;144;131;151m@[0m[38;2;144;135;154m@[0m[38;2;153;144;163m@[0m[38;2;154;145;164m@[0m[38;2;152;143;162m@[0m[38;2;151;142;161m@[0m[38;2;150;141;160m@[0m[38;2;150;141;160m@[0m[38;2;150;141;160m@[0m[38;2;150;141;162m@[0m[38;2;149;139;164m@[0m[38;2;148;138;163m@[0m[38;2;146;137;161m@[0m[38;2;146;136;161m@[0m[38;2;146;136;161m@[0m[38;2;146;137;158m@[0m[38;2;145;135;156m@[0m[38;2;144;134;155m@[0m[38;2;141;132;154m@[0m[38;2;141;131;156m@[0m[38;2;140;130;155m@[0m[38;2;139;129;154m@[0m[38;2;140;128;154m@[0m[38;2;140;128;153m@[0m[38;2;138;127;152m@[0m[38;2;135;126;151m@[0m[38;2;134;125;149m@[0m[38;2;131;125;150m@[0m[38;2;132;127;158m@[0m[38;2;133;127;163m@[0m[38;2;133;127;163m@[0m[38;2;99;95;121mB[0m[38;2;61;65;102mG[0m[38;2;66;73;121m#[0m[38;2;71;79;130m9[0m[38;2;76;87;136m9[0m[38;2;79;87;134m9[0m[38;2;79;85;131m9[0m[38;2;82;88;136mB[0m[38;2;89;95;138mB[0m[38;2;96;98;134mB[0m[38;2;122;117;155m@[0m[38;2;122;116;154m@[0m[38;2;102;97;130mB[0m[38;2;58;59;87mH[0m[38;2;56;47;69mh[0m[38;2;69;52;81mH[0m[38;2;72;52;81mH[0m[38;2;51;34;55m2[0m[38;2;41;27;47mX[0m[38;2;43;26;47mX[0m[38;2;47;33;54m2[0m[38;2;81;66;84mG[0m[38;2;90;68;88mS[0m[38;2;90;64;81mS[0m[38;2;58;39;53m5[0m[38;2;38;25;42ms[0m[38;2;55;42;61m3[0m[38;2;83;62;75mG[0m[38;2;49;31;45mA[0m[38;2;52;40;59m5[0m[38;2;84;62;76mG[0m[38;2;49;37;50m2[0m[38;2;31;31;47mX[0m[38;2;36;35;50mA[0m[38;2;35;32;46mX[0m[38;2;34;32;48mX[0m[38;2;30;30;44ms[0m");
	$display("[38;2;140;117;130m@[0m[38;2;140;116;130m@[0m[38;2;139;115;129m@[0m[38;2;138;115;129m@[0m[38;2;97;83;105m9[0m[38;2;88;67;85mS[0m[38;2;125;102;118m&[0m[38;2;80;66;89mS[0m[38;2;71;52;78mH[0m[38;2;77;56;78mH[0m[38;2;121;98;110mB[0m[38;2;101;85;104m9[0m[38;2;114;89;101mB[0m[38;2;140;113;127m@[0m[38;2;136;112;126m&[0m[38;2;130;106;120m&[0m[38;2;137;113;127m&[0m[38;2;141;117;130m@[0m[38;2;131;110;127m&[0m[38;2;83;67;89mS[0m[38;2;69;48;71mM[0m[38;2;72;52;73mM[0m[38;2;74;55;76mH[0m[38;2;66;48;70mM[0m[38;2;61;44;64m3[0m[38;2;57;43;61m3[0m[38;2;54;41;56m5[0m[38;2;51;39;51m2[0m[38;2;51;41;54m5[0m[38;2;62;53;74mM[0m[38;2;76;71;99mS[0m[38;2;84;84;119m9[0m[38;2;86;86;127m9[0m[38;2;86;87;128m9[0m[38;2;75;78;115m#[0m[38;2;66;69;101mS[0m[38;2;71;74;106mS[0m[38;2;72;75;109m#[0m[38;2;68;71;104mS[0m[38;2;62;67;97mG[0m[38;2;57;63;94mH[0m[38;2;57;60;87mH[0m[38;2;91;89;115m9[0m[38;2;144;142;167m@[0m[38;2;162;158;186m@[0m[38;2;158;154;183m@[0m[38;2;155;152;181m@[0m[38;2;148;145;175m@[0m[38;2;153;148;173m@[0m[38;2;157;148;168m@[0m[38;2;157;147;166m@[0m[38;2;156;147;166m@[0m[38;2;155;146;165m@[0m[38;2;154;145;164m@[0m[38;2;152;143;162m@[0m[38;2;150;141;160m@[0m[38;2;150;141;160m@[0m[38;2;150;141;160m@[0m[38;2;151;142;162m@[0m[38;2;150;141;162m@[0m[38;2;149;140;160m@[0m[38;2;148;139;160m@[0m[38;2;147;138;159m@[0m[38;2;148;137;161m@[0m[38;2;149;135;161m@[0m[38;2;148;135;158m@[0m[38;2;146;133;156m@[0m[38;2;146;132;157m@[0m[38;2;144;131;157m@[0m[38;2;144;130;156m@[0m[38;2;144;130;156m@[0m[38;2;142;129;154m@[0m[38;2;140;129;152m@[0m[38;2;138;128;150m@[0m[38;2;137;126;151m@[0m[38;2;136;126;150m@[0m[38;2;133;124;148m@[0m[38;2;132;123;149m@[0m[38;2;132;123;151m@[0m[38;2;132;125;158m@[0m[38;2;131;126;161m@[0m[38;2;131;125;161m@[0m[38;2;110;107;143m&[0m[38;2;80;84;126m9[0m[38;2;76;84;130m9[0m[38;2;89;98;139mB[0m[38;2;97;103;142m&[0m[38;2;101;106;145m&[0m[38;2;88;93;131mB[0m[38;2;76;81;119m9[0m[38;2;113;114;150m&[0m[38;2;123;117;155m@[0m[38;2;123;117;155m@[0m[38;2;101;96;130mB[0m[38;2;64;60;91mH[0m[38;2;70;51;82mH[0m[38;2;72;51;83mH[0m[38;2;72;52;81mH[0m[38;2;56;39;59m5[0m[38;2;40;27;44mX[0m[38;2;43;26;46mX[0m[38;2;46;32;53m2[0m[38;2;80;65;83mG[0m[38;2;89;67;86mS[0m[38;2;91;65;81mS[0m[38;2;62;41;54m3[0m[38;2;37;24;41ms[0m[38;2;48;36;56m2[0m[38;2;81;61;75mG[0m[38;2;51;30;45mA[0m[38;2;47;35;55m2[0m[38;2;82;63;78mG[0m[38;2;64;46;57m3[0m[38;2;31;31;44ms[0m[38;2;34;32;47mX[0m[38;2;34;31;47mX[0m[38;2;31;30;46ms[0m[38;2;29;29;43ms[0m");
	$display("[38;2;139;115;129m@[0m[38;2;140;116;130m@[0m[38;2;139;115;129m@[0m[38;2;138;114;128m@[0m[38;2;101;85;108m9[0m[38;2;74;58;78mH[0m[38;2;118;96;110mB[0m[38;2;85;71;92mS[0m[38;2;70;52;77mH[0m[38;2;70;51;74mM[0m[38;2;101;77;92m#[0m[38;2;114;95;111mB[0m[38;2;107;84;100m9[0m[38;2;138;112;126m&[0m[38;2;136;111;126m&[0m[38;2;133;109;123m&[0m[38;2;127;103;117m&[0m[38;2;138;114;128m@[0m[38;2;137;114;128m@[0m[38;2;98;82;101m9[0m[38;2;71;53;75mH[0m[38;2;88;67;92mS[0m[38;2;81;65;90mS[0m[38;2;56;46;62m3[0m[38;2;49;39;53m2[0m[38;2;50;38;52m2[0m[38;2;50;39;51m2[0m[38;2;61;54;72mM[0m[38;2;79;76;104m#[0m[38;2;86;86;125m9[0m[38;2;83;85;128m9[0m[38;2;87;88;129mB[0m[38;2;103;102;140m&[0m[38;2;90;92;126mB[0m[38;2;43;48;76m3[0m[38;2;60;63;93mG[0m[38;2;52;55;85mM[0m[38;2;43;47;75m3[0m[38;2;41;44;70m5[0m[38;2;45;47;71m3[0m[38;2;54;57;84mM[0m[38;2;64;65;95mG[0m[38;2;62;62;93mG[0m[38;2;68;69;95mG[0m[38;2;131;129;152m@[0m[38;2;161;158;185m@[0m[38;2;159;155;184m@[0m[38;2;157;154;183m@[0m[38;2;156;153;182m@[0m[38;2;153;149;173m@[0m[38;2;155;146;165m@[0m[38;2;156;146;165m@[0m[38;2;154;146;165m@[0m[38;2;153;144;163m@[0m[38;2;151;142;161m@[0m[38;2;150;142;161m@[0m[38;2;151;141;160m@[0m[38;2;151;141;160m@[0m[38;2;150;141;162m@[0m[38;2;150;141;162m@[0m[38;2;150;141;162m@[0m[38;2;149;139;160m@[0m[38;2;148;138;160m@[0m[38;2;149;137;159m@[0m[38;2;149;135;158m@[0m[38;2;149;135;158m@[0m[38;2;146;133;156m@[0m[38;2;144;134;155m@[0m[38;2;144;132;155m@[0m[38;2;145;131;157m@[0m[38;2;144;130;154m@[0m[38;2;143;129;153m@[0m[38;2;142;128;151m@[0m[38;2;141;127;150m@[0m[38;2;140;126;149m@[0m[38;2;138;125;149m@[0m[38;2;134;124;149m@[0m[38;2;132;123;148m@[0m[38;2;133;122;147m@[0m[38;2;133;121;147m@[0m[38;2;131;123;152m@[0m[38;2;131;125;158m@[0m[38;2;131;125;161m@[0m[38;2;123;117;152m@[0m[38;2;109;105;142m&[0m[38;2;98;100;136mB[0m[38;2;98;100;135mB[0m[38;2;101;101;137m&[0m[38;2;103;100;137m&[0m[38;2;117;113;150m@[0m[38;2;124;118;157m@[0m[38;2;124;117;156m@[0m[38;2;121;115;152m@[0m[38;2;91;82;114m9[0m[38;2;70;57;85mH[0m[38;2;67;50;79mM[0m[38;2;68;51;80mH[0m[38;2;70;50;80mH[0m[38;2;62;43;66mh[0m[38;2;43;29;45mX[0m[38;2;43;29;44mX[0m[38;2;44;30;48mA[0m[38;2;77;63;80mG[0m[38;2;89;67;85mS[0m[38;2;91;65;83mS[0m[38;2;63;43;56m3[0m[38;2;37;23;41ms[0m[38;2;43;31;49mA[0m[38;2;76;60;72mH[0m[38;2;50;32;42mA[0m[38;2;44;31;53mA[0m[38;2;79;63;79mG[0m[38;2;77;54;65mM[0m[38;2;36;29;42ms[0m[38;2;30;30;42ms[0m[38;2;33;32;45mX[0m[38;2;30;30;42ms[0m[38;2;28;28;39mr[0m");
	$display("[38;2;138;114;128m@[0m[38;2;139;115;129m@[0m[38;2;138;114;128m@[0m[38;2;137;113;128m&[0m[38;2;105;88;111mB[0m[38;2;67;54;75mM[0m[38;2;103;81;95m9[0m[38;2;90;74;94m#[0m[38;2;69;51;74mM[0m[38;2;70;51;74mM[0m[38;2;80;59;78mG[0m[38;2;116;94;111mB[0m[38;2;107;83;101m9[0m[38;2;136;110;123m&[0m[38;2;136;110;125m&[0m[38;2;137;110;125m&[0m[38;2;124;100;115m&[0m[38;2;126;103;117m&[0m[38;2;139;114;127m@[0m[38;2;117;98;116mB[0m[38;2;73;59;80mH[0m[38;2;73;59;81mH[0m[38;2;55;44;62m3[0m[38;2;50;38;52m2[0m[38;2;49;37;51m2[0m[38;2;54;44;57m5[0m[38;2;75;70;94mS[0m[38;2;87;85;125m9[0m[38;2;86;85;128m9[0m[38;2;94;93;132mB[0m[38;2;119;115;150m@[0m[38;2;144;141;170m@[0m[38;2;162;159;187m@[0m[38;2;110;112;138m&[0m[38;2;91;92;114m9[0m[38;2;112;113;137m&[0m[38;2;86;89;113m9[0m[38;2;49;51;77mh[0m[38;2;54;55;81mM[0m[38;2;79;81;108m#[0m[38;2;72;75;108m#[0m[38;2;71;76;109m#[0m[38;2;68;72;102mS[0m[38;2;60;64;93mG[0m[38;2;65;66;90mG[0m[38;2;146;142;167m@[0m[38;2;158;155;184m@[0m[38;2;156;153;182m@[0m[38;2;156;153;182m@[0m[38;2;155;152;179m@[0m[38;2;155;146;167m@[0m[38;2;155;146;164m@[0m[38;2;154;145;164m@[0m[38;2;153;144;163m@[0m[38;2;151;142;161m@[0m[38;2;152;142;161m@[0m[38;2;152;140;160m@[0m[38;2;154;141;161m@[0m[38;2;151;141;162m@[0m[38;2;152;139;162m@[0m[38;2;152;138;161m@[0m[38;2;152;138;161m@[0m[38;2;151;137;160m@[0m[38;2;150;136;159m@[0m[38;2;149;135;157m@[0m[38;2;149;135;158m@[0m[38;2;147;133;156m@[0m[38;2;146;132;156m@[0m[38;2;145;131;155m@[0m[38;2;145;131;157m@[0m[38;2;144;130;156m@[0m[38;2;142;128;154m@[0m[38;2;142;128;152m@[0m[38;2;141;127;149m@[0m[38;2;141;127;150m@[0m[38;2;139;126;150m@[0m[38;2;135;124;149m@[0m[38;2;133;122;148m@[0m[38;2;133;122;147m@[0m[38;2;134;120;146m@[0m[38;2;128;114;141m@[0m[38;2;113;103;131m&[0m[38;2;113;104;131m&[0m[38;2;114;107;133m&[0m[38;2;120;111;139m&[0m[38;2;121;112;141m&[0m[38;2;116;108;138m&[0m[38;2;112;105;136m&[0m[38;2;112;104;138m&[0m[38;2;111;105;138m&[0m[38;2;110;104;138m&[0m[38;2;106;100;134m&[0m[38;2;99;90;121mB[0m[38;2;85;71;95mS[0m[38;2;69;53;76mM[0m[38;2;65;45;75mM[0m[38;2;68;48;79mM[0m[38;2;68;48;79mM[0m[38;2;66;46;72mM[0m[38;2;48;33;49mA[0m[38;2;42;30;42mX[0m[38;2;40;29;46mX[0m[38;2;74;60;76mH[0m[38;2;90;66;84mS[0m[38;2;90;65;80mS[0m[38;2;66;46;58mh[0m[38;2;38;24;41ms[0m[38;2;40;27;47mX[0m[38;2;71;56;71mM[0m[38;2;50;32;43mA[0m[38;2;42;30;48mA[0m[38;2;76;61;77mH[0m[38;2;85;60;72mG[0m[38;2;43;32;44mA[0m[38;2;28;27;41mr[0m[38;2;33;31;45mX[0m[38;2;32;30;43ms[0m[38;2;26;24;36mi[0m");
	$display("[38;2;137;113;127m&[0m[38;2;137;113;127m&[0m[38;2;136;112;126m&[0m[38;2;136;112;126m&[0m[38;2;109;92;113mB[0m[38;2;66;54;75mM[0m[38;2;86;64;81mG[0m[38;2;91;72;93m#[0m[38;2;70;51;74mM[0m[38;2;69;49;71mM[0m[38;2;76;54;76mH[0m[38;2;113;87;107mB[0m[38;2;109;88;106mB[0m[38;2;133;107;120m&[0m[38;2;135;108;123m&[0m[38;2;136;108;123m&[0m[38;2;133;108;124m&[0m[38;2;111;88;104mB[0m[38;2;132;106;119m&[0m[38;2;134;109;124m&[0m[38;2;76;64;82mG[0m[38;2;48;37;51m2[0m[38;2;50;38;50m2[0m[38;2;49;37;50m2[0m[38;2;60;52;68mh[0m[38;2;82;79;110m#[0m[38;2;86;85;126m9[0m[38;2;94;93;130mB[0m[38;2;125;123;154m@[0m[38;2;153;150;179m@[0m[38;2;163;159;188m@[0m[38;2;163;158;187m@[0m[38;2;166;162;189m@[0m[38;2;149;150;176m@[0m[38;2;122;125;150m@[0m[38;2;97;101;128mB[0m[38;2;72;76;106m#[0m[38;2;84;91;128mB[0m[38;2;70;78;114m#[0m[38;2;66;74;106mS[0m[38;2;95;103;151m&[0m[38;2;92;101;150m&[0m[38;2;64;71;107mS[0m[38;2;84;91;130mB[0m[38;2;66;74;110mS[0m[38;2;116;116;141m&[0m[38;2;160;156;185m@[0m[38;2;156;153;182m@[0m[38;2;156;153;182m@[0m[38;2;154;152;180m@[0m[38;2;153;147;171m@[0m[38;2;155;145;164m@[0m[38;2;154;144;163m@[0m[38;2;153;143;162m@[0m[38;2;152;142;161m@[0m[38;2;154;141;161m@[0m[38;2;153;140;160m@[0m[38;2;153;140;161m@[0m[38;2;151;141;162m@[0m[38;2;151;140;162m@[0m[38;2;152;138;161m@[0m[38;2;152;138;161m@[0m[38;2;151;137;160m@[0m[38;2;150;136;158m@[0m[38;2;149;136;156m@[0m[38;2;148;134;156m@[0m[38;2;146;133;155m@[0m[38;2;146;132;157m@[0m[38;2;145;131;157m@[0m[38;2;145;131;157m@[0m[38;2;144;130;156m@[0m[38;2;143;129;154m@[0m[38;2;142;128;152m@[0m[38;2;141;127;149m@[0m[38;2;141;127;150m@[0m[38;2;140;126;150m@[0m[38;2;138;124;150m@[0m[38;2;136;122;148m@[0m[38;2;135;121;147m@[0m[38;2;134;120;146m@[0m[38;2;133;119;145m@[0m[38;2;124;114;139m&[0m[38;2;119;109;134m&[0m[38;2;116;104;131m&[0m[38;2;113;102;128m&[0m[38;2;117;104;129m&[0m[38;2;120;105;131m&[0m[38;2;119;103;129m&[0m[38;2;112;95;120mB[0m[38;2;104;86;112m9[0m[38;2;99;83;109m9[0m[38;2;100;84;110m9[0m[38;2;107;90;116mB[0m[38;2;117;98;125m&[0m[38;2;111;91;115mB[0m[38;2;78;56;84mG[0m[38;2;67;48;76mM[0m[38;2;69;49;77mM[0m[38;2;67;47;74mM[0m[38;2;58;39;59m3[0m[38;2;43;28;42mX[0m[38;2;39;27;45mX[0m[38;2;70;55;73mM[0m[38;2;89;66;80mS[0m[38;2;89;65;79mG[0m[38;2;72;49;62mh[0m[38;2;39;24;38ms[0m[38;2;40;26;46mX[0m[38;2;66;50;66mh[0m[38;2;51;33;44mA[0m[38;2;40;29;45mX[0m[38;2;73;59;75mH[0m[38;2;87;63;74mG[0m[38;2;53;38;48m2[0m[38;2;27;26;41mr[0m[38;2;30;29;45ms[0m[38;2;33;31;44mX[0m[38;2;26;24;36mi[0m");
	$display("[38;2;136;111;125m&[0m[38;2;136;111;125m&[0m[38;2;136;111;125m&[0m[38;2;137;112;125m&[0m[38;2;113;96;116mB[0m[38;2;69;54;78mH[0m[38;2;73;52;72mM[0m[38;2;80;61;83mG[0m[38;2;69;50;72mM[0m[38;2;68;48;70mM[0m[38;2;76;53;77mH[0m[38;2;106;80;106m9[0m[38;2;113;91;110mB[0m[38;2;130;104;117m&[0m[38;2;135;109;123m&[0m[38;2;134;108;123m&[0m[38;2;136;109;124m&[0m[38;2;122;99;114m&[0m[38;2;104;81;96m9[0m[38;2;137;110;123m&[0m[38;2;103;86;103m9[0m[38;2;53;41;58m5[0m[38;2;47;37;46mA[0m[38;2;63;58;74mM[0m[38;2;84;83;119m9[0m[38;2;86;86;126m9[0m[38;2;114;111;145m&[0m[38;2;151;148;176m@[0m[38;2;163;160;189m@[0m[38;2;161;158;188m@[0m[38;2;160;157;187m@[0m[38;2;160;157;187m@[0m[38;2;162;159;190m@[0m[38;2;137;141;171m@[0m[38;2;54;61;89mH[0m[38;2;53;57;86mM[0m[38;2;67;72;104mS[0m[38;2;87;98;139mB[0m[38;2;94;103;153m&[0m[38;2;88;99;147mB[0m[38;2;96;106;156m&[0m[38;2;97;108;157m&[0m[38;2;87;96;137mB[0m[38;2;116;124;163m@[0m[38;2;122;128;165m@[0m[38;2;134;134;162m@[0m[38;2;158;155;184m@[0m[38;2;156;153;182m@[0m[38;2;155;152;181m@[0m[38;2;154;152;178m@[0m[38;2;153;145;168m@[0m[38;2;157;144;163m@[0m[38;2;156;143;162m@[0m[38;2;157;144;163m@[0m[38;2;156;143;163m@[0m[38;2;154;141;161m@[0m[38;2;154;140;162m@[0m[38;2;154;140;163m@[0m[38;2;153;139;162m@[0m[38;2;153;139;162m@[0m[38;2;152;138;161m@[0m[38;2;152;138;161m@[0m[38;2;151;137;160m@[0m[38;2;149;136;158m@[0m[38;2;148;134;157m@[0m[38;2;146;133;153m@[0m[38;2;146;133;153m@[0m[38;2;146;132;155m@[0m[38;2;145;131;155m@[0m[38;2;145;131;157m@[0m[38;2;144;130;154m@[0m[38;2;143;129;152m@[0m[38;2;142;128;151m@[0m[38;2;140;126;149m@[0m[38;2;141;127;150m@[0m[38;2;141;127;150m@[0m[38;2;139;125;151m@[0m[38;2;137;123;149m@[0m[38;2;135;121;147m@[0m[38;2;134;120;146m@[0m[38;2;134;120;146m@[0m[38;2;129;119;144m@[0m[38;2;129;119;144m@[0m[38;2;127;117;142m@[0m[38;2;126;114;140m@[0m[38;2;127;113;139m@[0m[38;2;126;111;137m&[0m[38;2;125;109;136m&[0m[38;2;125;105;134m&[0m[38;2;124;104;132m&[0m[38;2;124;104;130m&[0m[38;2;122;101;127m&[0m[38;2;120;99;124m&[0m[38;2;118;98;124m&[0m[38;2;119;99;125m&[0m[38;2;107;86;110mB[0m[38;2;72;49;76mM[0m[38;2;66;45;74mM[0m[38;2;66;46;74mM[0m[38;2;63;44;65mh[0m[38;2;43;27;41mX[0m[38;2;39;25;44mX[0m[38;2;63;50;68mh[0m[38;2;88;65;80mG[0m[38;2;89;64;79mG[0m[38;2;78;55;67mH[0m[38;2;41;25;36ms[0m[38;2;38;25;41ms[0m[38;2;58;46;58m3[0m[38;2;50;33;44mA[0m[38;2;40;28;45mX[0m[38;2;65;52;66mh[0m[38;2;81;63;75mG[0m[38;2;63;46;55m3[0m[38;2;28;25;39mr[0m[38;2;29;27;42ms[0m[38;2;32;30;44ms[0m[38;2;26;24;36mi[0m");
	$display("[38;2;136;110;124m&[0m[38;2;136;110;124m&[0m[38;2;136;109;124m&[0m[38;2;138;110;124m&[0m[38;2;116;98;117mB[0m[38;2;70;56;78mH[0m[38;2;67;46;68mh[0m[38;2;68;49;71mM[0m[38;2;68;49;71mM[0m[38;2;67;48;70mM[0m[38;2;74;54;75mH[0m[38;2;101;78;105m9[0m[38;2;112;87;110mB[0m[38;2;129;105;117m&[0m[38;2;134;110;124m&[0m[38;2;133;109;123m&[0m[38;2;133;109;122m&[0m[38;2;135;110;123m&[0m[38;2;99;81;98m9[0m[38;2;109;85;98m9[0m[38;2;127;107;120m&[0m[38;2;68;57;74mH[0m[38;2;59;51;67mh[0m[38;2;87;85;118m9[0m[38;2;91;91;128mB[0m[38;2;131;128;157m@[0m[38;2;162;158;185m@[0m[38;2;161;158;187m@[0m[38;2;160;157;188m@[0m[38;2;160;157;188m@[0m[38;2;160;157;188m@[0m[38;2;160;157;188m@[0m[38;2;160;157;188m@[0m[38;2;161;159;189m@[0m[38;2;122;124;153m@[0m[38;2;79;83;117m9[0m[38;2;92;100;145m&[0m[38;2;82;91;133mB[0m[38;2;88;97;140mB[0m[38;2;108;119;158m@[0m[38;2;117;129;163m@[0m[38;2;122;134;167m@[0m[38;2;125;134;169m@[0m[38;2;117;126;163m@[0m[38;2;104;111;145m&[0m[38;2;151;147;175m@[0m[38;2;158;154;183m@[0m[38;2;156;152;182m@[0m[38;2;156;152;182m@[0m[38;2;152;149;172m@[0m[38;2;153;144;160m@[0m[38;2;158;146;161m@[0m[38;2;152;139;157m@[0m[38;2;130;115;139m@[0m[38;2;132;118;142m@[0m[38;2;153;140;161m@[0m[38;2;154;140;163m@[0m[38;2;153;139;162m@[0m[38;2;153;139;162m@[0m[38;2;153;139;162m@[0m[38;2;152;138;161m@[0m[38;2;151;137;160m@[0m[38;2;150;136;159m@[0m[38;2;149;136;157m@[0m[38;2;147;134;154m@[0m[38;2;146;133;153m@[0m[38;2;146;133;153m@[0m[38;2;146;132;155m@[0m[38;2;145;131;155m@[0m[38;2;145;131;155m@[0m[38;2;144;130;153m@[0m[38;2;142;128;151m@[0m[38;2;142;128;151m@[0m[38;2;141;127;150m@[0m[38;2;139;124;148m@[0m[38;2;129;114;139m@[0m[38;2;133;119;145m@[0m[38;2;137;123;149m@[0m[38;2;137;123;149m@[0m[38;2;136;122;146m@[0m[38;2;133;119;144m@[0m[38;2;128;118;143m@[0m[38;2;128;118;143m@[0m[38;2;125;116;141m@[0m[38;2;126;114;140m@[0m[38;2;127;113;139m@[0m[38;2;126;111;138m&[0m[38;2;125;109;136m&[0m[38;2;123;103;130m&[0m[38;2;120;100;127m&[0m[38;2;121;101;128m&[0m[38;2;119;99;126m&[0m[38;2;118;98;124m&[0m[38;2;117;97;123m&[0m[38;2;116;96;122mB[0m[38;2;117;96;120mB[0m[38;2;93;69;95m#[0m[38;2;68;45;73mM[0m[38;2;68;46;74mM[0m[38;2;64;44;65mh[0m[38;2;43;27;44mX[0m[38;2;39;26;43mX[0m[38;2;55;45;61m3[0m[38;2;87;65;80mG[0m[38;2;88;64;78mG[0m[38;2;84;58;71mH[0m[38;2;45;27;39mX[0m[38;2;36;24;39ms[0m[38;2;51;40;55m5[0m[38;2;48;31;44mA[0m[38;2;39;28;45mX[0m[38;2;58;45;56m3[0m[38;2;73;57;71mH[0m[38;2;74;53;63mM[0m[38;2;30;25;37mr[0m[38;2;27;26;39mr[0m[38;2;30;27;41ms[0m[38;2;27;26;36mr[0m");
	$display("[38;2;135;110;125m&[0m[38;2;136;110;125m&[0m[38;2;136;109;124m&[0m[38;2;137;110;124m&[0m[38;2;121;102;118m&[0m[38;2;72;59;81mH[0m[38;2;66;46;67mh[0m[38;2;67;48;70mM[0m[38;2;66;47;69mh[0m[38;2;65;46;69mh[0m[38;2;75;53;74mH[0m[38;2;100;77;106m9[0m[38;2;103;79;110m9[0m[38;2;124;99;114m&[0m[38;2;134;110;123m&[0m[38;2;133;109;122m&[0m[38;2;133;109;122m&[0m[38;2;136;109;122m&[0m[38;2;123;103;119m&[0m[38;2;79;63;80mG[0m[38;2;119;94;105mB[0m[38;2;104;88;102m9[0m[38;2;66;53;71mM[0m[38;2;83;76;107m#[0m[38;2;117;114;143m&[0m[38;2;164;161;185m@[0m[38;2;161;158;185m@[0m[38;2;160;157;186m@[0m[38;2;160;157;188m@[0m[38;2;160;157;188m@[0m[38;2;160;157;188m@[0m[38;2;160;157;188m@[0m[38;2;160;157;188m@[0m[38;2;160;157;188m@[0m[38;2;162;159;190m@[0m[38;2;145;144;175m@[0m[38;2;113;116;155m@[0m[38;2;97;105;150m&[0m[38;2;97;107;150m&[0m[38;2;114;123;157m@[0m[38;2;123;132;160m@[0m[38;2;131;137;164m@[0m[38;2;123;130;157m@[0m[38;2;117;120;152m@[0m[38;2;145;141;173m@[0m[38;2;159;154;184m@[0m[38;2;153;149;177m@[0m[38;2;150;144;170m@[0m[38;2;146;141;167m@[0m[38;2;140;132;152m@[0m[38;2;151;139;157m@[0m[38;2;135;121;143m@[0m[38;2;101;86;114m9[0m[38;2;111;95;123mB[0m[38;2;138;124;146m@[0m[38;2;154;141;163m@[0m[38;2;154;140;163m@[0m[38;2;153;139;162m@[0m[38;2;153;139;162m@[0m[38;2;153;139;162m@[0m[38;2;152;138;161m@[0m[38;2;151;137;160m@[0m[38;2;150;136;159m@[0m[38;2;149;136;157m@[0m[38;2;147;134;154m@[0m[38;2;146;133;153m@[0m[38;2;146;133;153m@[0m[38;2;146;132;155m@[0m[38;2;145;131;154m@[0m[38;2;145;131;154m@[0m[38;2;144;130;153m@[0m[38;2;142;128;151m@[0m[38;2;142;128;151m@[0m[38;2;140;126;149m@[0m[38;2;140;125;150m@[0m[38;2;127;111;137m&[0m[38;2;109;91;119mB[0m[38;2;105;88;116mB[0m[38;2;114;97;125m&[0m[38;2;123;107;134m&[0m[38;2;127;115;139m@[0m[38;2;128;118;143m@[0m[38;2;128;118;143m@[0m[38;2;125;116;141m@[0m[38;2;126;114;140m@[0m[38;2;127;113;139m@[0m[38;2;126;111;138m&[0m[38;2;125;109;136m&[0m[38;2;124;105;131m&[0m[38;2;121;101;127m&[0m[38;2;119;99;123m&[0m[38;2;119;99;125m&[0m[38;2;119;99;127m&[0m[38;2;117;97;125m&[0m[38;2;117;97;125m&[0m[38;2;117;95;121mB[0m[38;2;111;90;114mB[0m[38;2;76;53;77mH[0m[38;2;68;45;74mM[0m[38;2;65;43;65mh[0m[38;2;47;30;47mA[0m[38;2;40;27;43mX[0m[38;2;48;37;53m2[0m[38;2;84;64;78mG[0m[38;2;88;63;77mG[0m[38;2;87;61;74mG[0m[38;2;50;30;43mA[0m[38;2;36;22;39mr[0m[38;2;48;33;50m2[0m[38;2;46;30;42mX[0m[38;2;39;27;44mX[0m[38;2;56;40;53m5[0m[38;2;59;46;60m3[0m[38;2;80;59;71mH[0m[38;2;36;27;36ms[0m[38;2;25;23;37mi[0m[38;2;27;25;39mr[0m[38;2;28;27;37mr[0m");
	$display("[38;2;134;109;123m&[0m[38;2;134;109;123m&[0m[38;2;134;109;123m&[0m[38;2;135;110;123m&[0m[38;2;127;105;121m&[0m[38;2;78;64;85mG[0m[38;2;63;46;66mh[0m[38;2;67;47;69mh[0m[38;2;66;47;69mh[0m[38;2;65;46;68mh[0m[38;2;76;54;77mH[0m[38;2;99;76;107m9[0m[38;2;103;80;113m9[0m[38;2;120;97;113mB[0m[38;2;134;110;122m&[0m[38;2;133;109;122m&[0m[38;2;133;109;122m&[0m[38;2;133;108;121m&[0m[38;2;133;110;123m&[0m[38;2;100;84;101m9[0m[38;2;78;56;72mH[0m[38;2;124;99;108mB[0m[38;2;84;67;82mG[0m[38;2;77;60;75mH[0m[38;2;89;78;98m#[0m[38;2;132;126;147m@[0m[38;2;161;157;182m@[0m[38;2;162;158;188m@[0m[38;2;160;157;188m@[0m[38;2;160;157;187m@[0m[38;2;160;157;188m@[0m[38;2;159;157;188m@[0m[38;2;159;156;187m@[0m[38;2;159;156;187m@[0m[38;2;159;156;187m@[0m[38;2;161;158;188m@[0m[38;2;160;156;186m@[0m[38;2;151;149;178m@[0m[38;2;140;140;171m@[0m[38;2;133;134;165m@[0m[38;2;134;134;164m@[0m[38;2;140;138;168m@[0m[38;2;149;146;177m@[0m[38;2;157;152;182m@[0m[38;2;147;141;169m@[0m[38;2;138;130;155m@[0m[38;2;142;130;152m@[0m[38;2;150;136;156m@[0m[38;2;153;140;159m@[0m[38;2;147;133;153m@[0m[38;2;125;110;135m&[0m[38;2;113;97;122mB[0m[38;2;137;121;145m@[0m[38;2;155;142;159m@[0m[38;2;155;142;159m@[0m[38;2;154;141;159m@[0m[38;2;153;139;161m@[0m[38;2;153;139;162m@[0m[38;2;153;139;162m@[0m[38;2;152;138;161m@[0m[38;2;152;138;161m@[0m[38;2;151;137;160m@[0m[38;2;150;136;159m@[0m[38;2;149;135;156m@[0m[38;2;147;134;154m@[0m[38;2;146;133;153m@[0m[38;2;146;133;153m@[0m[38;2;146;132;155m@[0m[38;2;145;131;154m@[0m[38;2;145;131;154m@[0m[38;2;144;130;153m@[0m[38;2;142;128;151m@[0m[38;2;142;128;151m@[0m[38;2;141;127;150m@[0m[38;2;140;126;150m@[0m[38;2;140;126;151m@[0m[38;2;136;121;148m@[0m[38;2;121;105;131m&[0m[38;2;103;84;112m9[0m[38;2;95;73;104m#[0m[38;2;93;75;106m#[0m[38;2;118;108;135m&[0m[38;2;129;119;144m@[0m[38;2;126;117;142m@[0m[38;2;126;114;140m@[0m[38;2;127;113;139m@[0m[38;2;126;111;137m&[0m[38;2;126;109;137m&[0m[38;2;128;108;136m&[0m[38;2;125;105;133m&[0m[38;2;120;100;127m&[0m[38;2;120;100;127m&[0m[38;2;120;100;128m&[0m[38;2;118;98;126m&[0m[38;2;117;97;125m&[0m[38;2;116;96;123m&[0m[38;2;116;96;122mB[0m[38;2;94;73;94m#[0m[38;2;67;44;71mh[0m[38;2;65;43;64mh[0m[38;2;53;36;54m5[0m[38;2;47;33;49mA[0m[38;2;43;31;48mA[0m[38;2;78;61;78mG[0m[38;2;87;65;78mG[0m[38;2;86;64;76mG[0m[38;2;56;36;48m2[0m[38;2;36;21;38mr[0m[38;2;41;27;42mX[0m[38;2;40;25;40ms[0m[38;2;38;26;43ms[0m[38;2;56;41;54m5[0m[38;2;44;33;49mA[0m[38;2;78;60;74mH[0m[38;2;45;32;40mX[0m[38;2;24;23;35mi[0m[38;2;26;23;38mr[0m[38;2;26;25;35mi[0m");
	$display("[38;2;133;109;122m&[0m[38;2;133;109;122m&[0m[38;2;133;109;122m&[0m[38;2;134;109;122m&[0m[38;2;130;107;122m&[0m[38;2;87;72;92mS[0m[38;2;63;46;67mh[0m[38;2;66;47;67mh[0m[38;2;66;47;68mh[0m[38;2;65;46;68mh[0m[38;2;77;57;79mH[0m[38;2;101;77;105m9[0m[38;2;116;94;121mB[0m[38;2;130;111;130m&[0m[38;2;131;107;120m&[0m[38;2;132;108;121m&[0m[38;2;131;107;120m&[0m[38;2;131;107;120m&[0m[38;2;132;107;120m&[0m[38;2;126;105;118m&[0m[38;2;74;59;76mH[0m[38;2;86;63;75mG[0m[38;2;114;94;107mB[0m[38;2;75;56;75mH[0m[38;2;91;68;88mS[0m[38;2;106;91;108mB[0m[38;2;128;119;134m@[0m[38;2;145;140;162m@[0m[38;2;155;152;179m@[0m[38;2;160;157;187m@[0m[38;2;162;158;189m@[0m[38;2;161;157;188m@[0m[38;2;160;158;187m@[0m[38;2;160;157;187m@[0m[38;2;160;157;187m@[0m[38;2;159;157;186m@[0m[38;2;160;157;186m@[0m[38;2;160;157;186m@[0m[38;2;162;158;187m@[0m[38;2;161;158;187m@[0m[38;2;161;157;187m@[0m[38;2;155;151;178m@[0m[38;2;135;129;156m@[0m[38;2;125;115;137m&[0m[38;2;139;124;143m@[0m[38;2;153;135;153m@[0m[38;2;156;138;158m@[0m[38;2;155;137;158m@[0m[38;2;154;137;159m@[0m[38;2;151;134;156m@[0m[38;2;153;135;157m@[0m[38;2;156;139;160m@[0m[38;2;156;140;160m@[0m[38;2;153;139;158m@[0m[38;2;153;139;158m@[0m[38;2;151;138;157m@[0m[38;2;151;138;159m@[0m[38;2;153;139;161m@[0m[38;2;152;138;162m@[0m[38;2;152;138;161m@[0m[38;2;151;137;160m@[0m[38;2;150;136;159m@[0m[38;2;150;136;159m@[0m[38;2;148;134;156m@[0m[38;2;146;133;153m@[0m[38;2;146;133;153m@[0m[38;2;146;133;153m@[0m[38;2;146;132;155m@[0m[38;2;145;131;154m@[0m[38;2;144;130;153m@[0m[38;2;143;129;152m@[0m[38;2;142;128;151m@[0m[38;2;141;127;150m@[0m[38;2;141;127;150m@[0m[38;2;140;126;152m@[0m[38;2;139;125;151m@[0m[38;2;138;124;150m@[0m[38;2;138;124;148m@[0m[38;2;135;121;144m@[0m[38;2;127;111;136m&[0m[38;2;116;101;128m&[0m[38;2;122;111;138m&[0m[38;2;129;119;143m@[0m[38;2;127;118;143m@[0m[38;2;127;115;141m@[0m[38;2;127;113;139m@[0m[38;2;127;112;138m&[0m[38;2;125;110;137m&[0m[38;2;126;109;136m&[0m[38;2;125;107;135m&[0m[38;2;122;105;132m&[0m[38;2;122;103;131m&[0m[38;2;121;101;129m&[0m[38;2;120;100;128m&[0m[38;2;118;98;126m&[0m[38;2;117;97;125m&[0m[38;2;117;96;125m&[0m[38;2;111;90;111mB[0m[38;2;75;51;76mH[0m[38;2;65;43;65mh[0m[38;2;55;36;57m5[0m[38;2;54;38;56m5[0m[38;2;39;26;42ms[0m[38;2;69;54;71mM[0m[38;2;89;69;81mS[0m[38;2;86;65;77mG[0m[38;2;65;41;51m3[0m[38;2;36;21;36mr[0m[38;2;37;23;38ms[0m[38;2;37;22;39ms[0m[38;2;38;25;44ms[0m[38;2;58;43;58m3[0m[38;2;39;25;39ms[0m[38;2;68;53;68mM[0m[38;2;61;42;50m5[0m[38;2;22;20;33m;[0m[38;2;24;23;36mi[0m[38;2;21;21;32m;[0m");
	$display("[38;2;133;109;122m&[0m[38;2;133;109;122m&[0m[38;2;133;109;122m&[0m[38;2;133;109;122m&[0m[38;2;133;108;123m&[0m[38;2;97;81;100m9[0m[38;2;63;47;69mh[0m[38;2;64;46;65mh[0m[38;2;65;47;67mh[0m[38;2;63;47;68mh[0m[38;2;80;59;81mG[0m[38;2;99;78;104m9[0m[38;2;125;106;128m&[0m[38;2;140;125;142m@[0m[38;2;130;106;119m&[0m[38;2;131;107;120m&[0m[38;2;131;107;120m&[0m[38;2;131;107;120m&[0m[38;2;130;106;119m&[0m[38;2;131;107;120m&[0m[38;2;105;87;102m9[0m[38;2;61;45;62m3[0m[38;2;97;72;87m#[0m[38;2;101;81;98m9[0m[38;2;77;57;79mH[0m[38;2;125;104;126m&[0m[38;2;153;141;157m@[0m[38;2;142;133;149m@[0m[38;2;133;124;145m@[0m[38;2;136;127;152m@[0m[38;2;140;131;159m@[0m[38;2;145;136;168m@[0m[38;2;148;140;172m@[0m[38;2;151;146;174m@[0m[38;2;154;149;176m@[0m[38;2;155;149;179m@[0m[38;2;154;149;179m@[0m[38;2;150;146;174m@[0m[38;2;144;141;169m@[0m[38;2;134;130;156m@[0m[38;2;123;117;140m@[0m[38;2;116;106;125m&[0m[38;2;131;116;133m@[0m[38;2;152;133;152m@[0m[38;2;156;137;156m@[0m[38;2;155;136;155m@[0m[38;2;155;136;155m@[0m[38;2;154;135;155m@[0m[38;2;154;135;155m@[0m[38;2;154;134;155m@[0m[38;2;154;135;155m@[0m[38;2;154;135;157m@[0m[38;2;153;135;158m@[0m[38;2;152;137;158m@[0m[38;2;151;136;157m@[0m[38;2;150;137;157m@[0m[38;2;150;137;157m@[0m[38;2;151;138;158m@[0m[38;2;150;137;158m@[0m[38;2;151;138;159m@[0m[38;2;150;136;159m@[0m[38;2;150;136;158m@[0m[38;2;149;136;157m@[0m[38;2;147;134;155m@[0m[38;2;146;133;153m@[0m[38;2;146;133;153m@[0m[38;2;146;133;153m@[0m[38;2;146;132;155m@[0m[38;2;145;131;154m@[0m[38;2;144;130;153m@[0m[38;2;143;129;152m@[0m[38;2;142;128;151m@[0m[38;2;141;127;150m@[0m[38;2;140;126;149m@[0m[38;2;140;126;152m@[0m[38;2;139;125;151m@[0m[38;2;137;123;149m@[0m[38;2;136;122;146m@[0m[38;2;135;121;144m@[0m[38;2;135;121;144m@[0m[38;2;132;118;140m@[0m[38;2;107;100;121mB[0m[38;2;126;117;142m@[0m[38;2;128;118;143m@[0m[38;2;127;115;141m@[0m[38;2;127;113;139m@[0m[38;2;127;113;139m@[0m[38;2;125;111;137m&[0m[38;2;122;110;136m&[0m[38;2;123;109;135m&[0m[38;2;124;108;135m&[0m[38;2;122;105;132m&[0m[38;2;121;104;131m&[0m[38;2;121;102;130m&[0m[38;2;120;100;128m&[0m[38;2;118;98;126m&[0m[38;2;117;97;125m&[0m[38;2;118;98;122m&[0m[38;2;84;64;86mS[0m[38;2;62;42;64m3[0m[38;2;56;37;61m5[0m[38;2;62;41;63m3[0m[38;2;39;25;42ms[0m[38;2;57;42;59m3[0m[38;2;87;68;80mS[0m[38;2;89;67;79mS[0m[38;2;73;48;59mh[0m[38;2;38;21;36mr[0m[38;2;36;23;38mr[0m[38;2;37;22;38mr[0m[38;2;37;24;42ms[0m[38;2;59;44;59m3[0m[38;2;39;24;37ms[0m[38;2;51;38;54m5[0m[38;2;72;53;64mM[0m[38;2;27;24;35mi[0m[38;2;24;24;36mi[0m[38;2;23;22;33mi[0m");
	$display("[38;2;131;105;115m&[0m[38;2;132;108;121m&[0m[38;2;132;108;121m&[0m[38;2;132;107;120m&[0m[38;2;133;108;121m&[0m[38;2;108;92;109mB[0m[38;2;65;50;73mM[0m[38;2;64;45;64mh[0m[38;2;64;45;65mh[0m[38;2;63;46;65mh[0m[38;2;81;60;83mG[0m[38;2;100;77;106m9[0m[38;2;134;114;134m@[0m[38;2;145;134;150m@[0m[38;2;129;106;120m&[0m[38;2;131;107;120m&[0m[38;2;130;106;119m&[0m[38;2;130;106;119m&[0m[38;2;124;101;114m&[0m[38;2;124;99;112m&[0m[38;2;127;103;117m&[0m[38;2;77;59;80mG[0m[38;2;63;42;62m3[0m[38;2;109;84;96m9[0m[38;2;88;71;88mS[0m[38;2;81;62;84mG[0m[38;2;139;119;139m@[0m[38;2;164;146;165m@[0m[38;2;161;142;164m@[0m[38;2;156;137;159m@[0m[38;2;148;131;154m@[0m[38;2;121;106;130m&[0m[38;2;121;103;129m&[0m[38;2;126;110;137m&[0m[38;2;109;94;121mB[0m[38;2;120;103;130m&[0m[38;2;124;106;134m&[0m[38;2;121;105;131m&[0m[38;2;124;107;131m&[0m[38;2;132;114;134m@[0m[38;2;144;125;144m@[0m[38;2;153;135;153m@[0m[38;2;156;137;156m@[0m[38;2;154;135;154m@[0m[38;2;154;134;153m@[0m[38;2;155;134;153m@[0m[38;2;153;134;153m@[0m[38;2;153;134;153m@[0m[38;2;152;133;152m@[0m[38;2;151;132;151m@[0m[38;2;152;133;152m@[0m[38;2;152;134;153m@[0m[38;2;153;134;154m@[0m[38;2;154;135;157m@[0m[38;2;152;136;157m@[0m[38;2;150;136;156m@[0m[38;2;149;136;156m@[0m[38;2;149;136;156m@[0m[38;2;149;136;154m@[0m[38;2;151;138;155m@[0m[38;2;150;137;158m@[0m[38;2;150;137;158m@[0m[38;2;149;135;157m@[0m[38;2;147;134;155m@[0m[38;2;146;133;153m@[0m[38;2;146;133;153m@[0m[38;2;146;133;153m@[0m[38;2;146;132;155m@[0m[38;2;145;131;154m@[0m[38;2;144;130;153m@[0m[38;2;143;129;152m@[0m[38;2;141;127;150m@[0m[38;2;141;127;149m@[0m[38;2;141;128;150m@[0m[38;2;140;126;152m@[0m[38;2;139;125;151m@[0m[38;2;137;123;149m@[0m[38;2;136;122;146m@[0m[38;2;135;121;144m@[0m[38;2;135;121;144m@[0m[38;2;131;117;140m@[0m[38;2;120;109;133m&[0m[38;2;130;118;143m@[0m[38;2;127;118;143m@[0m[38;2;127;115;141m@[0m[38;2;127;113;139m@[0m[38;2;127;113;139m@[0m[38;2;125;111;137m&[0m[38;2;121;111;136m&[0m[38;2;121;110;135m&[0m[38;2;121;109;135m&[0m[38;2;121;108;134m&[0m[38;2;121;106;133m&[0m[38;2;120;105;131m&[0m[38;2;120;104;130m&[0m[38;2;119;102;129m&[0m[38;2;118;100;128m&[0m[38;2;120;100;127m&[0m[38;2;96;76;98m#[0m[38;2;65;43;67mh[0m[38;2;55;40;63m3[0m[38;2;63;45;68mh[0m[38;2;40;26;44mX[0m[38;2;43;30;47mA[0m[38;2;79;62;77mG[0m[38;2;91;69;81mS[0m[38;2;79;54;66mH[0m[38;2;41;23;38ms[0m[38;2;36;22;37mr[0m[38;2;37;23;38ms[0m[38;2;36;23;40ms[0m[38;2;58;43;58m3[0m[38;2;39;24;37ms[0m[38;2;38;25;42ms[0m[38;2;70;53;67mM[0m[38;2;44;31;40mX[0m[38;2;23;23;35mi[0m[38;2;22;21;33m;[0m");
	$display("[38;2;125;95;103mB[0m[38;2;134;106;120m&[0m[38;2;131;107;120m&[0m[38;2;131;107;120m&[0m[38;2;132;108;121m&[0m[38;2;119;100;116m&[0m[38;2;71;58;76mH[0m[38;2;62;43;62m3[0m[38;2;63;44;63mh[0m[38;2;63;44;63mh[0m[38;2;74;51;72mM[0m[38;2;98;73;99m#[0m[38;2;143;123;142m@[0m[38;2;149;139;155m@[0m[38;2;128;106;122m&[0m[38;2;131;106;119m&[0m[38;2;131;106;119m&[0m[38;2;132;106;119m&[0m[38;2;118;95;109mB[0m[38;2;114;90;102mB[0m[38;2;132;106;116m&[0m[38;2;103;86;99m9[0m[38;2;59;43;62m3[0m[38;2;85;60;80mG[0m[38;2;112;90;106mB[0m[38;2;79;61;78mG[0m[38;2;92;69;91mS[0m[38;2;147;126;144m@[0m[38;2;160;141;160m@[0m[38;2;158;139;159m@[0m[38;2;158;140;159m@[0m[38;2;151;134;152m@[0m[38;2;157;142;158m@[0m[38;2;157;142;159m@[0m[38;2;142;124;142m@[0m[38;2;155;134;152m@[0m[38;2;157;136;155m@[0m[38;2;158;137;155m@[0m[38;2;158;137;155m@[0m[38;2;157;137;156m@[0m[38;2;155;136;155m@[0m[38;2;153;134;153m@[0m[38;2;154;135;154m@[0m[38;2;153;134;153m@[0m[38;2;154;134;153m@[0m[38;2;155;134;153m@[0m[38;2;154;133;152m@[0m[38;2;153;133;152m@[0m[38;2;154;133;152m@[0m[38;2;153;132;151m@[0m[38;2;152;131;150m@[0m[38;2;151;132;151m@[0m[38;2;151;133;152m@[0m[38;2;151;134;156m@[0m[38;2;151;135;157m@[0m[38;2;151;136;157m@[0m[38;2;150;136;156m@[0m[38;2;149;136;156m@[0m[38;2;150;137;154m@[0m[38;2;150;137;154m@[0m[38;2;150;137;157m@[0m[38;2;150;137;157m@[0m[38;2;148;135;156m@[0m[38;2;147;134;154m@[0m[38;2;146;133;153m@[0m[38;2;146;132;155m@[0m[38;2;146;132;155m@[0m[38;2;146;132;155m@[0m[38;2;145;131;154m@[0m[38;2;144;130;153m@[0m[38;2;143;129;152m@[0m[38;2;141;127;150m@[0m[38;2;141;127;148m@[0m[38;2;141;128;148m@[0m[38;2;140;126;149m@[0m[38;2;139;125;149m@[0m[38;2;137;123;149m@[0m[38;2;136;122;146m@[0m[38;2;135;121;144m@[0m[38;2;135;121;144m@[0m[38;2;132;118;141m@[0m[38;2;133;118;142m@[0m[38;2;132;118;142m@[0m[38;2;130;117;143m@[0m[38;2;129;115;141m@[0m[38;2;128;114;140m@[0m[38;2;127;113;139m@[0m[38;2;125;111;137m&[0m[38;2;122;112;137m&[0m[38;2;121;111;136m&[0m[38;2;120;110;135m&[0m[38;2;120;110;135m&[0m[38;2;119;108;134m&[0m[38;2;119;106;132m&[0m[38;2;119;105;131m&[0m[38;2;116;104;130m&[0m[38;2;115;103;129m&[0m[38;2;118;103;129m&[0m[38;2;104;86;109m9[0m[38;2;66;45;69mh[0m[38;2;56;41;63m3[0m[38;2;63;46;69mh[0m[38;2;41;27;42mX[0m[38;2;38;25;41ms[0m[38;2;65;51;66mh[0m[38;2;88;69;81mS[0m[38;2;85;62;73mG[0m[38;2;46;27;41mX[0m[38;2;36;22;37mr[0m[38;2;37;23;38ms[0m[38;2;36;21;36mr[0m[38;2;57;44;56m3[0m[38;2;38;26;37ms[0m[38;2;31;21;37mr[0m[38;2;52;41;55m5[0m[38;2;60;44;53m3[0m[38;2;23;21;33mi[0m[38;2;19;20;31m;[0m");
	$display("[38;2;106;77;85m#[0m[38;2;133;103;115m&[0m[38;2;133;107;121m&[0m[38;2;133;107;120m&[0m[38;2;133;107;120m&[0m[38;2;127;105;117m&[0m[38;2;82;69;87mS[0m[38;2;61;43;62m3[0m[38;2;62;43;62m3[0m[38;2;63;44;62m3[0m[38;2;69;50;70mM[0m[38;2;85;62;84mG[0m[38;2;142;124;139m@[0m[38;2;153;144;160m@[0m[38;2;128;110;125m&[0m[38;2;130;106;119m&[0m[38;2;131;104;118m&[0m[38;2;130;105;116m&[0m[38;2;110;90;102m9[0m[38;2;102;80;93m#[0m[38;2;132;106;114m&[0m[38;2;125;102;114m&[0m[38;2;74;57;77mH[0m[38;2;71;49;68mM[0m[38;2;101;77;98m9[0m[38;2;109;88;103m9[0m[38;2;73;57;73mH[0m[38;2;100;77;97m#[0m[38;2;151;127;147m@[0m[38;2;157;139;157m@[0m[38;2;157;138;157m@[0m[38;2;155;136;155m@[0m[38;2;155;137;156m@[0m[38;2;156;137;155m@[0m[38;2;157;135;154m@[0m[38;2;156;135;154m@[0m[38;2;156;135;154m@[0m[38;2;155;134;153m@[0m[38;2;155;135;154m@[0m[38;2;154;135;154m@[0m[38;2;154;135;154m@[0m[38;2;153;134;153m@[0m[38;2;153;134;153m@[0m[38;2;153;134;153m@[0m[38;2;154;133;152m@[0m[38;2;154;133;152m@[0m[38;2;154;133;152m@[0m[38;2;154;133;152m@[0m[38;2;152;132;151m@[0m[38;2;151;132;151m@[0m[38;2;151;132;151m@[0m[38;2;152;133;152m@[0m[38;2;153;134;154m@[0m[38;2;152;134;156m@[0m[38;2;152;135;155m@[0m[38;2;151;136;154m@[0m[38;2;150;137;154m@[0m[38;2;150;137;154m@[0m[38;2;150;137;154m@[0m[38;2;150;137;154m@[0m[38;2;149;136;154m@[0m[38;2;149;136;154m@[0m[38;2;148;135;155m@[0m[38;2;146;133;153m@[0m[38;2;146;133;153m@[0m[38;2;146;132;155m@[0m[38;2;146;132;155m@[0m[38;2;146;132;155m@[0m[38;2;145;131;154m@[0m[38;2;144;130;153m@[0m[38;2;142;128;151m@[0m[38;2;141;127;150m@[0m[38;2;141;127;148m@[0m[38;2;141;128;148m@[0m[38;2;140;126;149m@[0m[38;2;139;125;149m@[0m[38;2;137;123;149m@[0m[38;2;136;122;148m@[0m[38;2;135;121;147m@[0m[38;2;135;121;145m@[0m[38;2;134;120;143m@[0m[38;2;132;118;143m@[0m[38;2;132;118;143m@[0m[38;2;131;117;143m@[0m[38;2;129;115;141m@[0m[38;2;128;114;140m@[0m[38;2;127;113;139m@[0m[38;2;127;113;139m@[0m[38;2;123;112;137m&[0m[38;2;120;111;136m&[0m[38;2;120;110;135m&[0m[38;2;120;110;135m&[0m[38;2;119;109;134m&[0m[38;2;120;107;133m&[0m[38;2;119;106;131m&[0m[38;2;116;106;131m&[0m[38;2;114;104;129m&[0m[38;2;115;104;130m&[0m[38;2;107;92;114mB[0m[38;2;68;47;71mM[0m[38;2;56;41;64m3[0m[38;2;63;47;69mh[0m[38;2;40;26;40ms[0m[38;2;36;23;38mr[0m[38;2;51;38;52m2[0m[38;2;83;66;81mG[0m[38;2;88;68;77mG[0m[38;2;55;33;44m2[0m[38;2;35;21;36mr[0m[38;2;37;23;39ms[0m[38;2;35;21;37mr[0m[38;2;55;42;54m5[0m[38;2;41;32;39mX[0m[38;2;25;20;34mi[0m[38;2;37;27;43ms[0m[38;2;65;50;62mh[0m[38;2;33;23;35mr[0m[38;2;20;19;29m;[0m");
	$display("[38;2;83;57;70mH[0m[38;2;124;97;105mB[0m[38;2;132;106;119m&[0m[38;2;131;105;118m&[0m[38;2;132;106;118m&[0m[38;2;130;106;115m&[0m[38;2;97;83;99m9[0m[38;2;60;46;64mh[0m[38;2;60;43;61m3[0m[38;2;61;42;61m3[0m[38;2;78;58;80mG[0m[38;2;100;77;103m9[0m[38;2;137;120;134m@[0m[38;2;152;144;159m@[0m[38;2;129;111;127m&[0m[38;2;125;102;114m&[0m[38;2;125;99;113m&[0m[38;2;131;104;114m&[0m[38;2;106;87;100m9[0m[38;2;89;67;81mS[0m[38;2;131;105;114m&[0m[38;2;131;106;115m&[0m[38;2;100;81;96m9[0m[38;2;59;43;61m3[0m[38;2;89;68;91mS[0m[38;2;102;79;102m9[0m[38;2;107;87;98m9[0m[38;2;73;53;72mM[0m[38;2;107;77;100m9[0m[38;2;152;127;146m@[0m[38;2;157;136;155m@[0m[38;2;154;134;153m@[0m[38;2;156;136;155m@[0m[38;2;155;135;154m@[0m[38;2;155;134;153m@[0m[38;2;156;135;154m@[0m[38;2;155;134;153m@[0m[38;2;154;133;152m@[0m[38;2;155;135;154m@[0m[38;2;155;135;154m@[0m[38;2;154;133;152m@[0m[38;2;155;135;154m@[0m[38;2;154;133;152m@[0m[38;2;154;133;152m@[0m[38;2;154;133;152m@[0m[38;2;154;133;152m@[0m[38;2;153;132;151m@[0m[38;2;153;133;152m@[0m[38;2;151;133;152m@[0m[38;2;152;133;152m@[0m[38;2;153;134;153m@[0m[38;2;153;134;155m@[0m[38;2;153;134;155m@[0m[38;2;153;134;156m@[0m[38;2;152;134;156m@[0m[38;2;150;135;156m@[0m[38;2;149;136;154m@[0m[38;2;150;137;154m@[0m[38;2;150;137;154m@[0m[38;2;150;137;154m@[0m[38;2;150;137;154m@[0m[38;2;149;136;153m@[0m[38;2;148;135;152m@[0m[38;2;146;133;152m@[0m[38;2;146;133;153m@[0m[38;2;146;132;155m@[0m[38;2;146;132;155m@[0m[38;2;146;132;155m@[0m[38;2;145;131;154m@[0m[38;2;144;130;153m@[0m[38;2;143;129;152m@[0m[38;2;141;127;150m@[0m[38;2;141;127;148m@[0m[38;2;141;128;148m@[0m[38;2;140;126;149m@[0m[38;2;139;125;149m@[0m[38;2;138;124;150m@[0m[38;2;137;123;147m@[0m[38;2;135;121;144m@[0m[38;2;135;121;144m@[0m[38;2;133;119;142m@[0m[38;2;133;119;142m@[0m[38;2;132;118;141m@[0m[38;2;131;117;143m@[0m[38;2;130;116;142m@[0m[38;2;128;114;140m@[0m[38;2;127;113;139m@[0m[38;2;125;112;138m&[0m[38;2;122;111;136m&[0m[38;2;120;111;136m&[0m[38;2;120;110;135m&[0m[38;2;120;110;135m&[0m[38;2;120;110;135m&[0m[38;2;118;108;133m&[0m[38;2;117;107;132m&[0m[38;2;116;106;131m&[0m[38;2;115;105;129m&[0m[38;2;115;105;130m&[0m[38;2;107;92;115mB[0m[38;2;69;48;72mM[0m[38;2;56;41;64m3[0m[38;2;60;44;66mh[0m[38;2;39;24;41ms[0m[38;2;37;23;39ms[0m[38;2;40;27;44mX[0m[38;2;75;59;75mH[0m[38;2;89;69;81mS[0m[38;2;64;43;54m3[0m[38;2;35;20;34mr[0m[38;2;37;23;38ms[0m[38;2;35;21;36mr[0m[38;2;51;38;52m2[0m[38;2;49;38;45m2[0m[38;2;21;19;32m;[0m[38;2;27;21;36mi[0m[38;2;50;40;54m5[0m[38;2;50;36;46m2[0m[38;2;18;18;30m:[0m");
	$display("[38;2;66;45;61mh[0m[38;2;108;80;88m9[0m[38;2;131;104;114m&[0m[38;2;130;104;115m&[0m[38;2;130;104;117m&[0m[38;2;131;105;116m&[0m[38;2;114;94;109mB[0m[38;2;65;51;71mM[0m[38;2;58;42;62m3[0m[38;2;62;42;61m3[0m[38;2;77;55;76mH[0m[38;2;104;81;106m9[0m[38;2;151;134;148m@[0m[38;2;155;147;165m@[0m[38;2;129;113;131m&[0m[38;2;122;96;109mB[0m[38;2;119;95;108mB[0m[38;2;133;105;115m&[0m[38;2;103;84;98m9[0m[38;2;76;54;71mH[0m[38;2;127;100;110m&[0m[38;2;131;107;116m&[0m[38;2;119;99;109mB[0m[38;2;68;51;68mM[0m[38;2;78;55;76mH[0m[38;2;100;74;102m9[0m[38;2;104;78;101m9[0m[38;2;104;83;98m9[0m[38;2;73;52;72mM[0m[38;2;107;80;101m9[0m[38;2;152;126;145m@[0m[38;2;157;136;154m@[0m[38;2;156;135;155m@[0m[38;2;156;135;154m@[0m[38;2;155;134;153m@[0m[38;2;154;133;152m@[0m[38;2;155;134;153m@[0m[38;2;155;134;153m@[0m[38;2;154;133;152m@[0m[38;2;155;134;153m@[0m[38;2;154;133;152m@[0m[38;2;155;134;153m@[0m[38;2;154;133;152m@[0m[38;2;154;133;152m@[0m[38;2;155;134;153m@[0m[38;2;155;134;153m@[0m[38;2;154;133;152m@[0m[38;2;153;133;152m@[0m[38;2;153;134;153m@[0m[38;2;153;134;155m@[0m[38;2;153;134;156m@[0m[38;2;153;134;156m@[0m[38;2;153;134;156m@[0m[38;2;153;134;156m@[0m[38;2;152;134;156m@[0m[38;2;150;135;156m@[0m[38;2;150;136;156m@[0m[38;2;149;136;156m@[0m[38;2;150;137;154m@[0m[38;2;150;137;154m@[0m[38;2;149;136;153m@[0m[38;2;149;136;153m@[0m[38;2;147;134;151m@[0m[38;2;146;133;152m@[0m[38;2;146;133;153m@[0m[38;2;146;132;155m@[0m[38;2;146;132;155m@[0m[38;2;146;132;155m@[0m[38;2;145;131;154m@[0m[38;2;144;130;153m@[0m[38;2;143;129;152m@[0m[38;2;141;127;150m@[0m[38;2;141;127;148m@[0m[38;2;141;128;148m@[0m[38;2;140;126;149m@[0m[38;2;139;125;148m@[0m[38;2;137;123;146m@[0m[38;2;136;122;145m@[0m[38;2;135;121;144m@[0m[38;2;135;121;144m@[0m[38;2;133;119;142m@[0m[38;2;132;118;141m@[0m[38;2;132;118;141m@[0m[38;2;131;117;143m@[0m[38;2;130;116;142m@[0m[38;2;128;114;140m@[0m[38;2;127;113;139m@[0m[38;2;125;112;138m&[0m[38;2;123;112;137m&[0m[38;2;120;111;136m&[0m[38;2;120;110;135m&[0m[38;2;120;110;135m&[0m[38;2;120;110;135m&[0m[38;2;118;108;133m&[0m[38;2;117;107;132m&[0m[38;2;116;106;131m&[0m[38;2;115;105;129m&[0m[38;2;115;105;130m&[0m[38;2;106;91;114mB[0m[38;2;68;48;72mM[0m[38;2;55;40;63m3[0m[38;2;53;38;55m5[0m[38;2;37;22;37mr[0m[38;2;37;23;38ms[0m[38;2;36;22;39mr[0m[38;2;62;48;63mh[0m[38;2;88;70;82mS[0m[38;2;75;53;64mM[0m[38;2;39;21;35mr[0m[38;2;36;22;37mr[0m[38;2;34;21;35mr[0m[38;2;44;32;48mA[0m[38;2;58;43;51m5[0m[38;2;23;20;32m;[0m[38;2;23;21;33mi[0m[38;2;33;26;41ms[0m[38;2;58;44;55m3[0m[38;2;28;21;30mi[0m");
	$display("[38;2;61;43;61m3[0m[38;2;85;59;70mH[0m[38;2;128;99;108m&[0m[38;2;130;104;117m&[0m[38;2;130;104;117m&[0m[38;2;130;104;117m&[0m[38;2;125;101;115m&[0m[38;2;78;64;81mG[0m[38;2;59;42;60m3[0m[38;2;60;41;60m3[0m[38;2;73;53;72mM[0m[38;2;103;79;104m9[0m[38;2;150;133;148m@[0m[38;2;157;149;166m@[0m[38;2;130;117;133m@[0m[38;2;116;92;106mB[0m[38;2;115;89;103mB[0m[38;2;132;104;114m&[0m[38;2;103;84;98m9[0m[38;2;64;45;62mh[0m[38;2;118;89;98mB[0m[38;2;133;107;117m&[0m[38;2;129;104;113m&[0m[38;2;88;71;86mS[0m[38;2;63;43;61m3[0m[38;2;97;71;95m#[0m[38;2;99;72;101m#[0m[38;2;120;95;112mB[0m[38;2;105;85;97m9[0m[38;2;72;53;72mM[0m[38;2;107;79;102m9[0m[38;2;153;126;145m@[0m[38;2;156;135;153m@[0m[38;2;156;135;154m@[0m[38;2;155;133;153m@[0m[38;2;154;133;152m@[0m[38;2;156;135;154m@[0m[38;2;155;134;153m@[0m[38;2;154;133;152m@[0m[38;2;156;135;154m@[0m[38;2;155;134;153m@[0m[38;2;155;134;153m@[0m[38;2;154;133;152m@[0m[38;2;154;133;152m@[0m[38;2;155;134;153m@[0m[38;2;155;134;153m@[0m[38;2;155;134;153m@[0m[38;2;154;134;153m@[0m[38;2;153;134;154m@[0m[38;2;153;134;155m@[0m[38;2;153;134;156m@[0m[38;2;153;134;156m@[0m[38;2;152;135;156m@[0m[38;2;151;136;157m@[0m[38;2;150;136;156m@[0m[38;2;149;136;156m@[0m[38;2;150;137;156m@[0m[38;2;149;136;156m@[0m[38;2;150;137;154m@[0m[38;2;150;137;154m@[0m[38;2;149;136;153m@[0m[38;2;149;136;153m@[0m[38;2;149;136;153m@[0m[38;2;147;134;151m@[0m[38;2;147;134;151m@[0m[38;2;147;133;155m@[0m[38;2;146;132;155m@[0m[38;2;146;132;155m@[0m[38;2;145;131;154m@[0m[38;2;144;130;153m@[0m[38;2;143;129;152m@[0m[38;2;141;127;150m@[0m[38;2;141;128;148m@[0m[38;2;141;128;148m@[0m[38;2;140;126;149m@[0m[38;2;139;125;148m@[0m[38;2;138;124;147m@[0m[38;2;137;123;147m@[0m[38;2;135;121;147m@[0m[38;2;135;121;144m@[0m[38;2;133;119;142m@[0m[38;2;132;118;143m@[0m[38;2;132;118;144m@[0m[38;2;132;118;144m@[0m[38;2;131;117;143m@[0m[38;2;129;115;141m@[0m[38;2;127;113;139m@[0m[38;2;126;112;138m&[0m[38;2;122;112;137m&[0m[38;2;121;111;136m&[0m[38;2;120;110;135m&[0m[38;2;120;110;135m&[0m[38;2;120;110;135m&[0m[38;2;119;109;134m&[0m[38;2;117;107;132m&[0m[38;2;117;106;132m&[0m[38;2;115;104;130m&[0m[38;2;115;105;130m&[0m[38;2;107;92;115mB[0m[38;2;70;49;74mM[0m[38;2;52;36;54m2[0m[38;2;42;28;44mX[0m[38;2;37;23;38ms[0m[38;2;36;22;37mr[0m[38;2;36;22;37mr[0m[38;2;48;35;50m2[0m[38;2;84;67;79mG[0m[38;2;82;60;67mH[0m[38;2;42;24;35ms[0m[38;2;36;21;37mr[0m[38;2;35;21;36mr[0m[38;2;39;26;42ms[0m[38;2;64;48;57m3[0m[38;2;27;21;31mi[0m[38;2;20;20;32m;[0m[38;2;25;19;33mi[0m[38;2;45;35;48mA[0m[38;2;45;33;40mX[0m");
	$display("[38;2;64;51;70mM[0m[38;2;66;46;60mh[0m[38;2;114;85;93m9[0m[38;2;131;104;115m&[0m[38;2;129;103;116m&[0m[38;2;129;103;116m&[0m[38;2;129;103;116m&[0m[38;2;96;80;97m#[0m[38;2;60;43;61m3[0m[38;2;59;40;58m3[0m[38;2;71;49;66mM[0m[38;2;102;76;102m9[0m[38;2;147;129;147m@[0m[38;2;157;150;166m@[0m[38;2;135;121;137m@[0m[38;2;111;89;104mB[0m[38;2;110;84;96m9[0m[38;2;131;103;112m&[0m[38;2;102;83;98m9[0m[38;2;56;41;58m5[0m[38;2;102;76;84m#[0m[38;2;132;107;114m&[0m[38;2;131;108;115m&[0m[38;2;109;89;103m9[0m[38;2;59;42;61m3[0m[38;2;83;58;81mG[0m[38;2;100;73;102m#[0m[38;2;131;105;127m&[0m[38;2;132;112;126m&[0m[38;2;102;83;95m9[0m[38;2;74;52;72mM[0m[38;2;111;83;103m9[0m[38;2;152;128;146m@[0m[38;2;156;135;155m@[0m[38;2;154;133;152m@[0m[38;2;156;135;154m@[0m[38;2;156;135;154m@[0m[38;2;154;133;152m@[0m[38;2;155;134;153m@[0m[38;2;155;134;153m@[0m[38;2;155;134;153m@[0m[38;2;155;134;153m@[0m[38;2;154;133;152m@[0m[38;2;155;134;153m@[0m[38;2;155;134;153m@[0m[38;2;155;134;153m@[0m[38;2;153;134;154m@[0m[38;2;153;134;154m@[0m[38;2;153;134;156m@[0m[38;2;153;134;156m@[0m[38;2;153;134;156m@[0m[38;2;151;136;157m@[0m[38;2;151;136;157m@[0m[38;2;150;137;157m@[0m[38;2;149;136;156m@[0m[38;2;149;136;156m@[0m[38;2;149;136;154m@[0m[38;2;150;137;154m@[0m[38;2;150;137;154m@[0m[38;2;149;136;153m@[0m[38;2;149;136;153m@[0m[38;2;149;136;153m@[0m[38;2;149;136;153m@[0m[38;2;148;135;152m@[0m[38;2;147;134;151m@[0m[38;2;145;132;152m@[0m[38;2;145;132;153m@[0m[38;2;145;131;154m@[0m[38;2;144;130;153m@[0m[38;2;143;129;152m@[0m[38;2;142;128;152m@[0m[38;2;141;127;150m@[0m[38;2;141;128;148m@[0m[38;2;141;127;148m@[0m[38;2;139;125;148m@[0m[38;2;139;124;148m@[0m[38;2;138;124;147m@[0m[38;2;137;123;147m@[0m[38;2;136;122;147m@[0m[38;2;136;121;145m@[0m[38;2;134;121;143m@[0m[38;2;133;120;143m@[0m[38;2;131;119;142m@[0m[38;2;123;110;131m&[0m[38;2;126;112;137m&[0m[38;2;130;115;142m@[0m[38;2;128;114;140m@[0m[38;2;126;112;137m&[0m[38;2;122;112;137m&[0m[38;2;121;111;136m&[0m[38;2;120;110;135m&[0m[38;2;120;110;135m&[0m[38;2;120;110;135m&[0m[38;2;118;108;133m&[0m[38;2;117;107;132m&[0m[38;2;120;106;132m&[0m[38;2;118;104;130m&[0m[38;2;116;105;131m&[0m[38;2;101;85;109m9[0m[38;2;70;50;76mM[0m[38;2;49;33;47mA[0m[38;2;36;22;37mr[0m[38;2;37;23;39ms[0m[38;2;36;22;37mr[0m[38;2;35;21;38mr[0m[38;2;39;26;42ms[0m[38;2;74;60;74mH[0m[38;2;85;64;71mG[0m[38;2;46;28;37mX[0m[38;2;35;21;37mr[0m[38;2;35;21;37mr[0m[38;2;35;22;39mr[0m[38;2;65;49;61mh[0m[38;2;38;26;36ms[0m[38;2;20;18;31m;[0m[38;2;22;18;30m;[0m[38;2;26;23;36mi[0m[38;2;46;38;48m2[0m");
	$display("[38;2;81;68;87mS[0m[38;2;58;42;62m3[0m[38;2;91;63;71mG[0m[38;2;127;99;107mB[0m[38;2;129;103;115m&[0m[38;2;129;103;116m&[0m[38;2;129;102;115m&[0m[38;2;114;94;106mB[0m[38;2;65;51;69mM[0m[38;2;57;37;56m5[0m[38;2;68;45;63mh[0m[38;2;96;71;97m#[0m[38;2;142;123;142m@[0m[38;2;159;152;166m@[0m[38;2;137;125;142m@[0m[38;2;108;88;106m9[0m[38;2;105;81;93m9[0m[38;2;130;103;111m&[0m[38;2;101;83;97m9[0m[38;2;55;38;58m5[0m[38;2;85;58;70mH[0m[38;2;127;100;107mB[0m[38;2;134;110;116m&[0m[38;2;126;100;112m&[0m[38;2;71;56;74mH[0m[38;2;66;45;63mh[0m[38;2;96;69;97m#[0m[38;2;120;96;117mB[0m[38;2;151;135;152m@[0m[38;2;126;107;120m&[0m[38;2;99;81;91m#[0m[38;2;74;51;72mM[0m[38;2;118;89;111mB[0m[38;2;157;131;152m@[0m[38;2;156;135;154m@[0m[38;2;156;135;154m@[0m[38;2;156;135;154m@[0m[38;2;153;132;151m@[0m[38;2;155;134;153m@[0m[38;2;155;134;153m@[0m[38;2;155;134;153m@[0m[38;2;155;134;153m@[0m[38;2;155;134;153m@[0m[38;2;154;134;153m@[0m[38;2;153;134;154m@[0m[38;2;153;134;155m@[0m[38;2;153;134;156m@[0m[38;2;153;134;156m@[0m[38;2;153;134;156m@[0m[38;2;153;135;157m@[0m[38;2;153;136;158m@[0m[38;2;152;137;158m@[0m[38;2;151;136;157m@[0m[38;2;150;137;157m@[0m[38;2;149;136;156m@[0m[38;2;149;136;156m@[0m[38;2;149;136;154m@[0m[38;2;150;137;154m@[0m[38;2;150;137;154m@[0m[38;2;149;136;153m@[0m[38;2;149;136;153m@[0m[38;2;149;136;153m@[0m[38;2;148;135;152m@[0m[38;2;147;134;151m@[0m[38;2;146;133;150m@[0m[38;2;144;131;150m@[0m[38;2;144;131;151m@[0m[38;2;145;131;154m@[0m[38;2;145;131;154m@[0m[38;2;144;130;153m@[0m[38;2;143;129;152m@[0m[38;2;142;128;150m@[0m[38;2;142;128;149m@[0m[38;2;142;129;148m@[0m[38;2;140;127;149m@[0m[38;2;139;125;149m@[0m[38;2;137;125;148m@[0m[38;2;135;124;147m@[0m[38;2;131;122;145m@[0m[38;2;126;118;139m@[0m[38;2;116;110;127m&[0m[38;2;100;93;111mB[0m[38;2;76;70;81mG[0m[38;2;39;31;40mX[0m[38;2;76;73;93mS[0m[38;2;129;118;143m@[0m[38;2;128;114;138m@[0m[38;2;127;113;136m&[0m[38;2;123;113;137m&[0m[38;2;121;111;136m&[0m[38;2;120;110;135m&[0m[38;2;120;110;135m&[0m[38;2;120;110;135m&[0m[38;2;119;109;134m&[0m[38;2;117;107;132m&[0m[38;2;118;105;131m&[0m[38;2;117;105;131m&[0m[38;2;115;103;125m&[0m[38;2;83;64;88mS[0m[38;2;65;45;69mh[0m[38;2;42;26;41mX[0m[38;2;36;23;37mr[0m[38;2;37;23;38ms[0m[38;2;37;23;38ms[0m[38;2;36;22;37mr[0m[38;2;36;22;38mr[0m[38;2;65;52;65mh[0m[38;2;88;66;76mG[0m[38;2;52;33;42mA[0m[38;2;34;21;36mr[0m[38;2;36;21;37mr[0m[38;2;35;21;38mr[0m[38;2;58;43;58m3[0m[38;2;53;36;46m2[0m[38;2;21;18;31m;[0m[38;2;22;20;33m;[0m[38;2;22;20;33m;[0m[38;2;26;24;36mi[0m");
	$display("[38;2;104;88;103m9[0m[38;2;62;49;68mh[0m[38;2;70;45;60mh[0m[38;2;117;86;93m9[0m[38;2;129;103;111m&[0m[38;2;128;102;115m&[0m[38;2;129;102;115m&[0m[38;2;124;101;111m&[0m[38;2;81;68;84mG[0m[38;2;55;39;57m5[0m[38;2;63;42;61m3[0m[38;2;89;67;91mS[0m[38;2;113;90;113mB[0m[38;2;146;130;146m@[0m[38;2;141;130;145m@[0m[38;2;110;90;109mB[0m[38;2;104;78;93m#[0m[38;2;128;101;108m&[0m[38;2;100;82;95m9[0m[38;2;56;38;56m5[0m[38;2;68;44;60mh[0m[38;2;117;92;98mB[0m[38;2;133;108;114m&[0m[38;2;131;106;116m&[0m[38;2;92;76;90m#[0m[38;2;56;37;56m5[0m[38;2;85;60;83mG[0m[38;2;112;87;108mB[0m[38;2;156;138;156m@[0m[38;2;144;132;149m@[0m[38;2;123;101;113m&[0m[38;2;90;70;86mS[0m[38;2;77;53;73mH[0m[38;2;127;98;121m&[0m[38;2;157;135;154m@[0m[38;2;155;135;154m@[0m[38;2;155;135;154m@[0m[38;2;154;133;152m@[0m[38;2;155;135;154m@[0m[38;2;153;136;155m@[0m[38;2;153;136;155m@[0m[38;2;153;135;155m@[0m[38;2;154;135;155m@[0m[38;2;154;135;155m@[0m[38;2;154;135;157m@[0m[38;2;154;135;157m@[0m[38;2;153;135;157m@[0m[38;2;153;136;157m@[0m[38;2;153;136;158m@[0m[38;2;152;137;157m@[0m[38;2;151;137;157m@[0m[38;2;150;137;157m@[0m[38;2;150;137;157m@[0m[38;2;150;137;157m@[0m[38;2;149;136;156m@[0m[38;2;149;136;156m@[0m[38;2;149;136;154m@[0m[38;2;150;137;154m@[0m[38;2;150;137;154m@[0m[38;2;149;136;153m@[0m[38;2;149;136;153m@[0m[38;2;149;136;153m@[0m[38;2;148;135;152m@[0m[38;2;147;134;151m@[0m[38;2;146;133;150m@[0m[38;2;143;130;150m@[0m[38;2;143;130;151m@[0m[38;2;144;131;153m@[0m[38;2;144;130;153m@[0m[38;2;145;131;153m@[0m[38;2;142;129;148m@[0m[38;2;137;126;144m@[0m[38;2;134;123;144m@[0m[38;2;130;119;140m@[0m[38;2;123;112;134m&[0m[38;2;116;105;126m&[0m[38;2;105;94;114mB[0m[38;2;94;80;101m#[0m[38;2;81;66;83mG[0m[38;2;70;53;68mM[0m[38;2;64;41;57m3[0m[38;2;49;28;42mA[0m[38;2;30;15;26m;[0m[38;2;15;7;18m [0m[38;2;52;50;69mh[0m[38;2;127;117;141m@[0m[38;2;128;115;138m@[0m[38;2;127;113;136m&[0m[38;2;123;112;137m&[0m[38;2;121;111;136m&[0m[38;2;120;110;135m&[0m[38;2;120;110;135m&[0m[38;2;120;110;135m&[0m[38;2;119;109;134m&[0m[38;2;117;107;132m&[0m[38;2;117;106;131m&[0m[38;2;118;106;131m&[0m[38;2;100;84;105m9[0m[38;2;69;50;74mM[0m[38;2;52;33;50m2[0m[38;2;39;22;37ms[0m[38;2;38;22;38ms[0m[38;2;37;23;38ms[0m[38;2;36;22;37mr[0m[38;2;36;22;37mr[0m[38;2;35;20;36mr[0m[38;2;57;44;58m3[0m[38;2;87;66;77mG[0m[38;2;58;37;46m2[0m[38;2;35;20;36mr[0m[38;2;36;22;37mr[0m[38;2;36;21;36mr[0m[38;2;49;35;50m2[0m[38;2;65;46;56m3[0m[38;2;24;20;32m;[0m[38;2;21;21;33m;[0m[38;2;22;19;33m;[0m[38;2;21;17;29m:[0m");
	$display("[38;2;120;97;109mB[0m[38;2;80;67;85mG[0m[38;2;56;40;57m5[0m[38;2;95;67;75mS[0m[38;2;127;100;107mB[0m[38;2;126;101;112m&[0m[38;2;127;101;112m&[0m[38;2;128;102;112m&[0m[38;2;104;85;98m9[0m[38;2;57;43;61m3[0m[38;2;60;40;57m3[0m[38;2;83;61;83mG[0m[38;2;92;69;98m#[0m[38;2;101;78;105m9[0m[38;2;126;104;124m&[0m[38;2;111;90;107mB[0m[38;2;101;77;95m#[0m[38;2;126;99;105mB[0m[38;2;99;81;95m#[0m[38;2;56;38;57m5[0m[38;2;58;37;53m5[0m[38;2;102;76;84m#[0m[38;2;130;104;112m&[0m[38;2;133;110;118m&[0m[38;2;111;92;103mB[0m[38;2;60;41;60m3[0m[38;2;71;47;67mM[0m[38;2;102;77;98m9[0m[38;2;150;131;147m@[0m[38;2;157;146;162m@[0m[38;2;135;125;140m@[0m[38;2;117;95;111mB[0m[38;2;77;56;74mH[0m[38;2;84;58;80mG[0m[38;2;134;111;131m&[0m[38;2;157;138;155m@[0m[38;2;155;136;155m@[0m[38;2;155;136;156m@[0m[38;2;155;136;157m@[0m[38;2;155;136;158m@[0m[38;2;155;136;158m@[0m[38;2;156;137;159m@[0m[38;2;155;137;158m@[0m[38;2;155;138;158m@[0m[38;2;154;137;157m@[0m[38;2;154;138;157m@[0m[38;2;153;139;158m@[0m[38;2;152;139;158m@[0m[38;2;151;139;159m@[0m[38;2;151;138;158m@[0m[38;2;150;137;157m@[0m[38;2;150;137;157m@[0m[38;2;150;137;157m@[0m[38;2;150;137;157m@[0m[38;2;149;136;156m@[0m[38;2;149;136;156m@[0m[38;2;149;136;154m@[0m[38;2;150;137;154m@[0m[38;2;150;137;154m@[0m[38;2;149;136;153m@[0m[38;2;149;136;153m@[0m[38;2;149;136;153m@[0m[38;2;148;135;152m@[0m[38;2;146;133;150m@[0m[38;2;145;132;149m@[0m[38;2;143;130;150m@[0m[38;2;142;129;149m@[0m[38;2;142;129;150m@[0m[38;2;144;130;149m@[0m[38;2;117;101;114mB[0m[38;2;75;54;67mM[0m[38;2;67;47;61mh[0m[38;2;68;48;61mh[0m[38;2;65;45;59m3[0m[38;2;66;42;57m3[0m[38;2;68;41;57m3[0m[38;2;71;42;58mh[0m[38;2;80;46;63mM[0m[38;2;90;54;70mH[0m[38;2;99;62;77mS[0m[38;2;107;67;83m#[0m[38;2;109;71;89m#[0m[38;2;94;65;83mS[0m[38;2;67;53;75mM[0m[38;2;94;88;113m9[0m[38;2;128;116;139m@[0m[38;2;129;114;137m@[0m[38;2;127;113;136m&[0m[38;2;122;112;137m&[0m[38;2;121;111;136m&[0m[38;2;120;110;135m&[0m[38;2;120;110;135m&[0m[38;2;120;110;135m&[0m[38;2;118;108;133m&[0m[38;2;117;107;132m&[0m[38;2;121;106;133m&[0m[38;2;113;96;119mB[0m[38;2;76;56;82mH[0m[38;2;54;36;56m5[0m[38;2;43;27;42mX[0m[38;2;39;23;37ms[0m[38;2;38;22;36mr[0m[38;2;37;23;36mr[0m[38;2;36;23;36mr[0m[38;2;36;22;37mr[0m[38;2;35;20;36mr[0m[38;2;52;40;56m5[0m[38;2;86;65;78mG[0m[38;2;63;40;51m5[0m[38;2;35;20;35mr[0m[38;2;36;21;37mr[0m[38;2;37;22;38mr[0m[38;2;39;27;44mX[0m[38;2;70;51;63mM[0m[38;2;32;24;34mr[0m[38;2;20;19;32m;[0m[38;2;22;18;32m;[0m[38;2;20;15;28m:[0m");
	$display("[38;2;106;81;97m9[0m[38;2;103;85;98m9[0m[38;2;60;46;63m3[0m[38;2;70;47;60mh[0m[38;2;117;89;96m9[0m[38;2;127;101;109m&[0m[38;2;126;100;109m&[0m[38;2;127;100;109m&[0m[38;2;119;96;108mB[0m[38;2;71;57;75mH[0m[38;2;55;36;56m5[0m[38;2;70;49;67mM[0m[38;2;91;68;93mS[0m[38;2;89;65;97mS[0m[38;2;91;66;92mS[0m[38;2;108;84;98m9[0m[38;2;95;72;91m#[0m[38;2;124;95;104mB[0m[38;2;101;81;96m9[0m[38;2;55;37;58m5[0m[38;2;54;35;53m2[0m[38;2;82;55;65mH[0m[38;2;126;97;105mB[0m[38;2;133;109;116m&[0m[38;2;125;102;110m&[0m[38;2;72;55;73mH[0m[38;2;59;38;57m5[0m[38;2;90;67;87mS[0m[38;2;137;120;133m@[0m[38;2;158;146;162m@[0m[38;2;154;144;160m@[0m[38;2;130;112;129m&[0m[38;2;107;85;98m9[0m[38;2;64;45;63mh[0m[38;2;94;69;91m#[0m[38;2;146;125;143m@[0m[38;2;156;140;158m@[0m[38;2;155;138;158m@[0m[38;2;155;139;158m@[0m[38;2;155;139;158m@[0m[38;2;155;139;158m@[0m[38;2;155;139;158m@[0m[38;2;154;140;158m@[0m[38;2;154;141;157m@[0m[38;2;154;141;157m@[0m[38;2;154;141;158m@[0m[38;2;154;141;158m@[0m[38;2;153;140;157m@[0m[38;2;152;139;158m@[0m[38;2;151;138;157m@[0m[38;2;150;137;157m@[0m[38;2;151;138;158m@[0m[38;2;150;137;157m@[0m[38;2;150;137;157m@[0m[38;2;149;136;156m@[0m[38;2;149;136;154m@[0m[38;2;150;137;154m@[0m[38;2;150;137;154m@[0m[38;2;150;137;154m@[0m[38;2;149;136;153m@[0m[38;2;149;136;153m@[0m[38;2;149;136;153m@[0m[38;2;148;135;152m@[0m[38;2;146;133;150m@[0m[38;2;144;131;148m@[0m[38;2;143;130;149m@[0m[38;2;142;129;149m@[0m[38;2;144;131;150m@[0m[38;2;101;85;101m9[0m[38;2;50;26;40mX[0m[38;2;62;34;49m5[0m[38;2;82;49;64mM[0m[38;2;96;59;76mG[0m[38;2;106;67;84m#[0m[38;2;112;72;88m#[0m[38;2;115;76;93m9[0m[38;2;118;79;97m9[0m[38;2;119;83;101mB[0m[38;2;119;87;107mB[0m[38;2;120;92;111mB[0m[38;2;122;99;120m&[0m[38;2;125;108;130m&[0m[38;2;129;115;139m@[0m[38;2;133;119;146m@[0m[38;2;134;119;144m@[0m[38;2;130;116;140m@[0m[38;2;128;114;138m@[0m[38;2;127;113;136m&[0m[38;2;123;112;137m&[0m[38;2;121;111;136m&[0m[38;2;120;110;135m&[0m[38;2;120;110;135m&[0m[38;2;120;110;135m&[0m[38;2;119;109;134m&[0m[38;2;117;108;133m&[0m[38;2;118;104;127m&[0m[38;2;86;65;89mS[0m[38;2;59;39;59m3[0m[38;2;40;24;38ms[0m[38;2;42;29;44mX[0m[38;2;38;24;39ms[0m[38;2;37;23;38ms[0m[38;2;37;23;36mr[0m[38;2;36;23;35mr[0m[38;2;36;22;37mr[0m[38;2;35;21;36mr[0m[38;2;52;37;55m5[0m[38;2;85;66;78mG[0m[38;2;66;43;57m3[0m[38;2;35;20;34mr[0m[38;2;35;22;37mr[0m[38;2;37;23;39ms[0m[38;2;35;22;38mr[0m[38;2;64;48;61mh[0m[38;2;47;34;43mA[0m[38;2;19;18;31m;[0m[38;2;21;19;32m;[0m[38;2;18;17;28m:[0m");
	$display("[38;2;93;70;96m#[0m[38;2;105;84;100m9[0m[38;2;79;63;80mG[0m[38;2;57;40;56m5[0m[38;2;97;69;77mS[0m[38;2;125;98;107mB[0m[38;2;124;98;107mB[0m[38;2;125;99;107mB[0m[38;2;125;99;108mB[0m[38;2;93;77;90m#[0m[38;2;52;40;58m5[0m[38;2;59;39;58m3[0m[38;2;81;58;79mG[0m[38;2;90;67;96mS[0m[38;2;92;68;97m#[0m[38;2;107;82;97m9[0m[38;2;92;69;89mS[0m[38;2;115;88;99m9[0m[38;2;105;84;98m9[0m[38;2;56;38;57m5[0m[38;2;54;35;53m2[0m[38;2;62;40;53m5[0m[38;2;114;84;91m9[0m[38;2;131;105;112m&[0m[38;2;131;108;114m&[0m[38;2;92;74;88m#[0m[38;2;53;34;52m2[0m[38;2;79;57;76mH[0m[38;2;120;101;118m&[0m[38;2;157;143;160m@[0m[38;2;157;144;161m@[0m[38;2;149;137;155m@[0m[38;2;123;103;116m&[0m[38;2;85;67;81mG[0m[38;2;65;43;64mh[0m[38;2;109;85;107m9[0m[38;2;153;137;154m@[0m[38;2;155;142;158m@[0m[38;2;154;141;158m@[0m[38;2;154;141;158m@[0m[38;2;154;141;158m@[0m[38;2;154;141;158m@[0m[38;2;154;141;158m@[0m[38;2;154;141;158m@[0m[38;2;154;141;158m@[0m[38;2;154;141;158m@[0m[38;2;154;141;158m@[0m[38;2;154;141;158m@[0m[38;2;151;138;157m@[0m[38;2;150;137;157m@[0m[38;2;150;137;157m@[0m[38;2;150;137;157m@[0m[38;2;149;136;156m@[0m[38;2;149;136;156m@[0m[38;2;149;136;155m@[0m[38;2;149;136;153m@[0m[38;2;150;137;154m@[0m[38;2;150;137;154m@[0m[38;2;149;136;153m@[0m[38;2;149;136;153m@[0m[38;2;149;136;153m@[0m[38;2;149;136;153m@[0m[38;2;148;135;152m@[0m[38;2;147;134;151m@[0m[38;2;145;132;149m@[0m[38;2;143;130;149m@[0m[38;2;143;130;150m@[0m[38;2;143;130;148m@[0m[38;2;112;99;118mB[0m[38;2;102;85;105m9[0m[38;2;122;100;119m&[0m[38;2;126;102;120m&[0m[38;2;128;103;124m&[0m[38;2;128;105;125m&[0m[38;2;128;108;129m&[0m[38;2;129;112;134m&[0m[38;2;131;117;139m@[0m[38;2;132;119;141m@[0m[38;2;134;121;144m@[0m[38;2;134;121;145m@[0m[38;2;134;121;145m@[0m[38;2;133;120;143m@[0m[38;2;133;119;142m@[0m[38;2;132;118;144m@[0m[38;2;131;117;143m@[0m[38;2;130;116;142m@[0m[38;2;128;114;138m@[0m[38;2;127;113;136m&[0m[38;2;122;112;136m&[0m[38;2;121;111;136m&[0m[38;2;120;110;135m&[0m[38;2;120;110;135m&[0m[38;2;120;110;135m&[0m[38;2;120;110;134m&[0m[38;2;120;107;129m&[0m[38;2;93;76;97m#[0m[38;2;62;42;64m3[0m[38;2;41;25;39ms[0m[38;2;38;23;36mr[0m[38;2;42;28;40mX[0m[38;2;39;25;37ms[0m[38;2;37;24;36mr[0m[38;2;37;23;38ms[0m[38;2;37;23;38ms[0m[38;2;37;23;39ms[0m[38;2;38;23;37ms[0m[38;2;53;40;56m5[0m[38;2;86;65;77mG[0m[38;2;69;45;58mh[0m[38;2;36;20;35mr[0m[38;2;35;22;37mr[0m[38;2;37;23;38ms[0m[38;2;35;22;37mr[0m[38;2;49;37;51m2[0m[38;2;64;47;55m3[0m[38;2;23;18;30m;[0m[38;2;20;20;33m;[0m[38;2;18;18;29m:[0m");
	$display("[38;2;75;54;74mH[0m[38;2;85;63;81mG[0m[38;2;91;72;86mS[0m[38;2;60;43;62m3[0m[38;2;75;48;59mh[0m[38;2;119;90;95mB[0m[38;2;125;99;108mB[0m[38;2;125;99;108mB[0m[38;2;125;98;107mB[0m[38;2;113;92;102mB[0m[38;2;64;51;67mh[0m[38;2;54;35;54m5[0m[38;2;68;47;62mh[0m[38;2;91;69;93mS[0m[38;2;94;69;99m#[0m[38;2;107;81;98m9[0m[38;2;94;72;93m#[0m[38;2;105;78;96m9[0m[38;2;106;87;99m9[0m[38;2;58;40;58m3[0m[38;2;56;35;53m5[0m[38;2;54;34;51m2[0m[38;2;92;64;72mG[0m[38;2;128;99;107mB[0m[38;2;133;109;114m&[0m[38;2;108;88;101m9[0m[38;2;55;39;57m5[0m[38;2;70;47;68mM[0m[38;2;105;81;103m9[0m[38;2;152;135;152m@[0m[38;2;157;144;161m@[0m[38;2;156;145;162m@[0m[38;2;137;124;140m@[0m[38;2;111;90;105mB[0m[38;2;62;43;62m3[0m[38;2;78;54;75mH[0m[38;2;131;110;129m&[0m[38;2;157;143;160m@[0m[38;2;154;141;158m@[0m[38;2;154;141;158m@[0m[38;2;154;141;158m@[0m[38;2;154;141;158m@[0m[38;2;154;141;158m@[0m[38;2;154;141;158m@[0m[38;2;154;141;158m@[0m[38;2;154;141;158m@[0m[38;2;153;140;157m@[0m[38;2;152;139;157m@[0m[38;2;150;137;157m@[0m[38;2;150;137;157m@[0m[38;2;150;137;157m@[0m[38;2;150;137;157m@[0m[38;2;149;136;156m@[0m[38;2;149;136;156m@[0m[38;2;149;136;155m@[0m[38;2;150;137;154m@[0m[38;2;150;137;154m@[0m[38;2;149;136;153m@[0m[38;2;149;136;153m@[0m[38;2;149;136;153m@[0m[38;2;149;136;153m@[0m[38;2;149;136;153m@[0m[38;2;147;134;151m@[0m[38;2;147;134;151m@[0m[38;2;145;132;149m@[0m[38;2;143;130;149m@[0m[38;2;143;130;150m@[0m[38;2;142;129;149m@[0m[38;2;145;131;151m@[0m[38;2;146;133;152m@[0m[38;2;143;131;150m@[0m[38;2;142;130;149m@[0m[38;2;142;130;150m@[0m[38;2;142;130;151m@[0m[38;2;142;128;152m@[0m[38;2;139;126;149m@[0m[38;2;139;125;148m@[0m[38;2;138;124;147m@[0m[38;2;136;122;145m@[0m[38;2;135;121;144m@[0m[38;2;134;120;143m@[0m[38;2;133;119;142m@[0m[38;2;132;118;141m@[0m[38;2;131;117;143m@[0m[38;2;131;117;143m@[0m[38;2;130;116;142m@[0m[38;2;129;115;138m@[0m[38;2;126;113;136m&[0m[38;2;122;111;136m&[0m[38;2;121;111;136m&[0m[38;2;120;110;135m&[0m[38;2;120;110;135m&[0m[38;2;120;110;135m&[0m[38;2;122;110;134m&[0m[38;2;104;86;106m9[0m[38;2;67;47;69mh[0m[38;2;45;27;44mX[0m[38;2;37;23;38ms[0m[38;2;37;23;38ms[0m[38;2;40;26;39ms[0m[38;2;41;28;39mX[0m[38;2;37;24;34mr[0m[38;2;37;23;37mr[0m[38;2;37;23;37mr[0m[38;2;38;27;42ms[0m[38;2;51;37;50m2[0m[38;2;57;45;60m3[0m[38;2;86;64;77mG[0m[38;2;71;47;60mh[0m[38;2;37;21;36mr[0m[38;2;35;22;37mr[0m[38;2;36;22;37mr[0m[38;2;36;22;38mr[0m[38;2;36;27;41ms[0m[38;2;67;52;63mh[0m[38;2;35;25;36mr[0m[38;2;19;19;32m;[0m[38;2;18;18;29m:[0m");
	$display("\033[31m \033[5m     //   / /     //   ) )     //   ) )     //   ) )     //   ) )\033[0m");
    $display("\033[31m \033[5m    //____       //___/ /     //___/ /     //   / /     //___/ /\033[0m");
    $display("\033[31m \033[5m   / ____       / ___ (      / ___ (      //   / /     / ___ (\033[0m");
    $display("\033[31m \033[5m  //           //   | |     //   | |     //   / /     //   | |\033[0m");
    $display("\033[31m \033[5m //____/ /    //    | |    //    | |    ((___/ /     //    | |\033[0m");
end endtask

task display_pass; begin
	$display("[38;2;178;138;79m&[0m[38;2;179;139;79m&[0m[38;2;179;139;80m&[0m[38;2;180;140;80m&[0m[38;2;180;140;80m&[0m[38;2;180;140;81m&[0m[38;2;180;140;81m&[0m[38;2;181;141;82m&[0m[38;2;181;141;82m&[0m[38;2;181;141;81m&[0m[38;2;183;143;82m&[0m[38;2;183;143;83m&[0m[38;2;182;142;82m&[0m[38;2;182;142;82m&[0m[38;2;183;143;83m&[0m[38;2;184;144;84m&[0m[38;2;184;144;82m&[0m[38;2;183;143;81m&[0m[38;2;183;143;83m&[0m[38;2;183;143;84m&[0m[38;2;183;143;84m&[0m[38;2;183;143;84m&[0m[38;2;184;144;85m&[0m[38;2;183;143;84m&[0m[38;2;183;143;84m&[0m[38;2;183;143;84m&[0m[38;2;184;144;85m&[0m[38;2;184;144;85m&[0m[38;2;184;144;83m&[0m[38;2;184;144;83m&[0m[38;2;184;144;83m&[0m[38;2;184;144;83m&[0m[38;2;184;144;83m&[0m[38;2;184;144;83m&[0m[38;2;184;144;83m&[0m[38;2;184;144;83m&[0m[38;2;184;144;83m&[0m[38;2;184;144;83m&[0m[38;2;183;143;82m&[0m[38;2;183;143;82m&[0m[38;2;184;144;83m&[0m[38;2;183;143;82m&[0m[38;2;183;143;83m&[0m[38;2;181;142;79m&[0m[38;2;181;137;78m&[0m[38;2;116;60;35mH[0m[38;2;75;7;6mX[0m[38;2;77;7;9mX[0m[38;2;70;9;7mX[0m[38;2;67;22;11mA[0m[38;2;89;60;41mM[0m[38;2;124;104;78m9[0m[38;2;169;150;116m@[0m[38;2;190;172;134m@[0m[38;2;192;174;136m@[0m[38;2;192;176;138m@[0m[38;2;192;177;136m@[0m[38;2;194;179;136m@[0m[38;2;201;186;146m@[0m[38;2;180;164;127m@[0m[38;2;186;170;134m@[0m[38;2;192;177;139m@[0m[38;2;196;181;142m@[0m[38;2;195;180;140m@[0m[38;2;196;181;141m@[0m[38;2;195;180;141m@[0m[38;2;195;180;141m@[0m[38;2;196;181;142m@[0m[38;2;194;179;140m@[0m[38;2;196;179;139m@[0m[38;2;196;178;138m@[0m[38;2;188;170;132m@[0m[38;2;164;145;112m&[0m[38;2;135;115;87mB[0m[38;2;94;74;52mH[0m[38;2;57;39;23m2[0m[38;2;47;22;13ms[0m[38;2;58;19;13mX[0m[38;2;74;17;13mA[0m[38;2;83;13;10mA[0m[38;2;91;12;11mA[0m[38;2;95;13;10m2[0m[38;2;92;14;9m2[0m[38;2;91;14;10m2[0m[38;2;89;10;12mA[0m[38;2;89;10;12mA[0m[38;2;85;14;6mA[0m[38;2;101;38;19m3[0m[38;2;148;93;61m9[0m[38;2;165;117;70mB[0m[38;2;159;117;63mB[0m[38;2;159;117;66mB[0m[38;2;159;118;66mB[0m[38;2;157;116;63mB[0m[38;2;156;115;64mB[0m[38;2;156;114;63mB[0m[38;2;157;115;65mB[0m[38;2;170;128;80m&[0m[38;2;171;129;81m&[0m[38;2;171;129;81m&[0m[38;2;172;130;82m&[0m[38;2;173;130;82m&[0m[38;2;148;111;66m9[0m[38;2;115;83;44mG[0m[38;2;135;94;56m#[0m[38;2;161;116;71mB[0m[38;2;177;137;87m&[0m[38;2;185;148;95m@[0m[38;2;187;152;95m@[0m[38;2;187;152;96m@[0m[38;2;188;151;96m@[0m[38;2;188;151;96m@[0m[38;2;188;151;96m@[0m[38;2;189;152;96m@[0m[38;2;187;150;95m@[0m[38;2;187;151;94m@[0m[38;2;187;151;92m@[0m[38;2;187;151;92m@[0m[38;2;188;151;96m@[0m[38;2;162;125;73mB[0m[38;2;143;104;57m9[0m[38;2;145;103;58m9[0m[38;2;146;103;59m9[0m[38;2;145;103;60m9[0m[38;2;143;100;58m9[0m[38;2;160;117;69mB[0m[38;2;177;138;79m&[0m[38;2;193;156;94m@[0m[38;2;194;157;99m@[0m[38;2;177;136;80m&[0m[38;2;183;141;87m&[0m[38;2;188;150;91m@[0m[38;2;186;152;87m&[0m[38;2;186;152;90m@[0m[38;2;185;149;87m&[0m");
	$display("[38;2;175;135;79m&[0m[38;2;176;136;80m&[0m[38;2;176;136;80m&[0m[38;2;177;137;81m&[0m[38;2;177;137;81m&[0m[38;2;177;138;80m&[0m[38;2;177;138;80m&[0m[38;2;178;138;81m&[0m[38;2;179;139;81m&[0m[38;2;178;139;80m&[0m[38;2;179;140;81m&[0m[38;2;180;140;82m&[0m[38;2;179;140;81m&[0m[38;2;179;140;81m&[0m[38;2;180;140;81m&[0m[38;2;181;141;81m&[0m[38;2;181;141;81m&[0m[38;2;181;141;80m&[0m[38;2;181;141;81m&[0m[38;2;181;141;83m&[0m[38;2;182;142;83m&[0m[38;2;182;142;83m&[0m[38;2;182;142;83m&[0m[38;2;182;142;83m&[0m[38;2;182;142;83m&[0m[38;2;182;142;83m&[0m[38;2;182;142;83m&[0m[38;2;182;142;82m&[0m[38;2;182;142;81m&[0m[38;2;182;142;81m&[0m[38;2;182;142;81m&[0m[38;2;182;142;81m&[0m[38;2;182;142;81m&[0m[38;2;182;142;81m&[0m[38;2;182;142;81m&[0m[38;2;182;142;81m&[0m[38;2;182;142;81m&[0m[38;2;181;141;80m&[0m[38;2;180;140;79m&[0m[38;2;181;141;80m&[0m[38;2;182;142;81m&[0m[38;2;181;140;79m&[0m[38;2;180;139;76m&[0m[38;2;181;140;77m&[0m[38;2;155;105;63m9[0m[38;2;81;17;8mA[0m[38;2;79;5;9mX[0m[38;2;71;4;4ms[0m[38;2;74;26;15m2[0m[38;2;125;97;72m#[0m[38;2;168;150;116m@[0m[38;2;182;164;127m@[0m[38;2;195;177;139m@[0m[38;2;186;168;130m@[0m[38;2;194;176;138m@[0m[38;2;192;175;139m@[0m[38;2;190;175;136m@[0m[38;2;208;193;154m@[0m[38;2;176;161;124m@[0m[38;2;181;165;131m@[0m[38;2;177;161;128m@[0m[38;2;190;175;138m@[0m[38;2;211;196;156m@[0m[38;2;195;180;142m@[0m[38;2;175;159;123m@[0m[38;2;189;174;136m@[0m[38;2;195;180;138m@[0m[38;2;201;186;146m@[0m[38;2;202;186;149m@[0m[38;2;193;177;138m@[0m[38;2;195;179;140m@[0m[38;2;204;188;150m@[0m[38;2;205;188;150m@[0m[38;2;189;173;134m@[0m[38;2;185;168;131m@[0m[38;2;167;151;116m@[0m[38;2;122;106;78m9[0m[38;2;77;57;38mh[0m[38;2;50;29;13mX[0m[38;2;50;20;9ms[0m[38;2;65;16;12mX[0m[38;2;78;12;10mA[0m[38;2;85;12;7mA[0m[38;2;84;11;5mA[0m[38;2;83;8;6mX[0m[38;2;83;8;9mA[0m[38;2;83;7;6mX[0m[38;2;82;8;5mX[0m[38;2;88;21;12m2[0m[38;2;132;76;48mS[0m[38;2;157;112;67mB[0m[38;2;155;115;64mB[0m[38;2;155;114;64mB[0m[38;2;155;113;64mB[0m[38;2;154;112;63m9[0m[38;2;153;111;63m9[0m[38;2;155;112;65mB[0m[38;2;170;128;80m&[0m[38;2;172;130;82m&[0m[38;2;173;131;83m&[0m[38;2;173;131;83m&[0m[38;2;174;131;84m&[0m[38;2;147;109;65m9[0m[38;2;113;80;42mG[0m[38;2;134;92;56m#[0m[38;2;160;115;71mB[0m[38;2;175;135;86m&[0m[38;2;186;149;96m@[0m[38;2;187;152;95m@[0m[38;2;186;151;94m@[0m[38;2;187;150;95m@[0m[38;2;186;151;96m@[0m[38;2;186;151;96m@[0m[38;2;186;151;96m@[0m[38;2;185;150;95m@[0m[38;2;186;149;94m@[0m[38;2;186;149;93m@[0m[38;2;186;149;93m@[0m[38;2;187;150;97m@[0m[38;2;162;125;74mB[0m[38;2;143;104;58m9[0m[38;2;145;103;58m9[0m[38;2;146;103;59m9[0m[38;2;145;103;60m9[0m[38;2;143;101;58m9[0m[38;2;155;113;66mB[0m[38;2;171;131;77m&[0m[38;2;186;149;91m&[0m[38;2;187;151;94m@[0m[38;2;167;128;74mB[0m[38;2;172;132;82m&[0m[38;2;183;144;92m&[0m[38;2;178;141;89m&[0m[38;2;150;113;72mB[0m[38;2;109;78;48mG[0m");
	$display("[38;2;173;134;80m&[0m[38;2;173;134;80m&[0m[38;2;173;134;80m&[0m[38;2;174;135;81m&[0m[38;2;174;135;80m&[0m[38;2;175;136;80m&[0m[38;2;176;137;81m&[0m[38;2;176;137;80m&[0m[38;2;176;138;80m&[0m[38;2;177;138;80m&[0m[38;2;177;138;81m&[0m[38;2;177;138;81m&[0m[38;2;177;138;81m&[0m[38;2;177;138;81m&[0m[38;2;178;137;81m&[0m[38;2;178;138;81m&[0m[38;2;178;138;81m&[0m[38;2;179;138;81m&[0m[38;2;179;139;81m&[0m[38;2;179;139;80m&[0m[38;2;179;139;80m&[0m[38;2;179;139;80m&[0m[38;2;179;139;80m&[0m[38;2;179;139;80m&[0m[38;2;180;140;80m&[0m[38;2;180;140;80m&[0m[38;2;180;140;80m&[0m[38;2;180;140;79m&[0m[38;2;180;140;79m&[0m[38;2;181;141;79m&[0m[38;2;180;140;79m&[0m[38;2;180;140;79m&[0m[38;2;180;140;79m&[0m[38;2;179;139;78m&[0m[38;2;179;139;78m&[0m[38;2;179;139;78m&[0m[38;2;180;140;79m&[0m[38;2;179;139;78m&[0m[38;2;179;139;78m&[0m[38;2;179;139;78m&[0m[38;2;178;138;77m&[0m[38;2;179;137;79m&[0m[38;2;178;137;77m&[0m[38;2;176;135;79m&[0m[38;2;122;66;41mG[0m[38;2;75;7;7mX[0m[38;2;70;2;3ms[0m[38;2;76;24;14mA[0m[38;2;162;130;105m&[0m[38;2;188;169;133m@[0m[38;2;168;152;112m@[0m[38;2;193;176;140m@[0m[38;2;183;167;130m@[0m[38;2;190;174;136m@[0m[38;2;192;176;137m@[0m[38;2;188;172;134m@[0m[38;2;208;192;157m@[0m[38;2;177;161;127m@[0m[38;2;145;129;94mB[0m[38;2;176;160;127m@[0m[38;2;178;163;129m@[0m[38;2;203;188;150m@[0m[38;2;216;199;160m@[0m[38;2;186;168;134m@[0m[38;2;123;105;74m9[0m[38;2;105;89;58mS[0m[38;2;183;168;132m@[0m[38;2;194;179;138m@[0m[38;2;211;195;160m@[0m[38;2;201;185;150m@[0m[38;2;171;155;120m@[0m[38;2;190;174;141m@[0m[38;2;205;189;153m@[0m[38;2;211;196;157m@[0m[38;2;192;176;135m@[0m[38;2;190;174;132m@[0m[38;2;196;180;139m@[0m[38;2;187;171;134m@[0m[38;2;154;139;107m&[0m[38;2;91;78;52mH[0m[38;2;47;31;15mX[0m[38;2;48;19;13ms[0m[38;2;59;14;13mX[0m[38;2;70;10;6mX[0m[38;2;76;7;5mX[0m[38;2;80;6;5mX[0m[38;2;81;8;6mX[0m[38;2;83;9;7mX[0m[38;2;81;7;4mX[0m[38;2;76;13;3mX[0m[38;2;120;70;46mG[0m[38;2;152;111;64m9[0m[38;2;153;112;61m9[0m[38;2;152;110;62m9[0m[38;2;152;110;62m9[0m[38;2;151;109;62m9[0m[38;2;153;110;64m9[0m[38;2;170;128;80m&[0m[38;2;173;131;83m&[0m[38;2;173;132;84m&[0m[38;2;173;132;84m&[0m[38;2;174;133;85m&[0m[38;2;146;109;66m9[0m[38;2;113;78;41mG[0m[38;2;131;92;55m#[0m[38;2;157;114;71mB[0m[38;2;174;133;84m&[0m[38;2;184;147;95m&[0m[38;2;185;151;95m@[0m[38;2;183;150;94m&[0m[38;2;185;149;96m@[0m[38;2;184;150;96m@[0m[38;2;184;150;96m@[0m[38;2;184;150;96m@[0m[38;2;184;149;95m@[0m[38;2;185;148;95m@[0m[38;2;185;148;94m&[0m[38;2;185;148;93m&[0m[38;2;186;149;96m@[0m[38;2;160;123;75mB[0m[38;2;140;101;57m#[0m[38;2;136;95;56m#[0m[38;2;130;89;54m#[0m[38;2;125;83;50mS[0m[38;2;121;79;47mS[0m[38;2;124;83;50mS[0m[38;2;130;90;55m#[0m[38;2;134;93;59m#[0m[38;2;135;95;62m#[0m[38;2;128;88;54m#[0m[38;2;124;87;54mS[0m[38;2;100;69;39mH[0m[38;2;79;53;32mh[0m[38;2;54;31;20mA[0m[38;2;39;23;12ms[0m");
	$display("[38;2;172;133;78m&[0m[38;2;173;134;79m&[0m[38;2;173;134;78m&[0m[38;2;173;134;79m&[0m[38;2;173;134;78m&[0m[38;2;174;135;78m&[0m[38;2;174;135;78m&[0m[38;2;174;135;76m&[0m[38;2;174;134;76m&[0m[38;2;173;135;77m&[0m[38;2;175;136;79m&[0m[38;2;174;136;79m&[0m[38;2;175;137;79m&[0m[38;2;176;137;80m&[0m[38;2;177;136;80m&[0m[38;2;177;136;80m&[0m[38;2;177;136;80m&[0m[38;2;177;136;80m&[0m[38;2;177;136;80m&[0m[38;2;177;136;81m&[0m[38;2;177;136;81m&[0m[38;2;177;136;81m&[0m[38;2;178;137;82m&[0m[38;2;178;137;80m&[0m[38;2;178;137;80m&[0m[38;2;177;137;79m&[0m[38;2;177;137;79m&[0m[38;2;178;137;79m&[0m[38;2;177;137;79m&[0m[38;2;178;137;79m&[0m[38;2;178;137;79m&[0m[38;2;178;137;79m&[0m[38;2;177;137;79m&[0m[38;2;176;136;78m&[0m[38;2;177;136;78m&[0m[38;2;177;137;78m&[0m[38;2;177;137;78m&[0m[38;2;177;136;78m&[0m[38;2;177;137;78m&[0m[38;2;177;137;78m&[0m[38;2;176;136;77m&[0m[38;2;176;134;78m&[0m[38;2;174;135;78m&[0m[38;2;173;129;82m&[0m[38;2;107;47;29mM[0m[38;2;68;2;3ms[0m[38;2;78;30;16m2[0m[38;2;178;145;120m@[0m[38;2;183;165;131m@[0m[38;2;145;132;93mB[0m[38;2;196;181;143m@[0m[38;2;179;163;128m@[0m[38;2;185;170;132m@[0m[38;2;194;179;140m@[0m[38;2;184;169;130m@[0m[38;2;197;182;145m@[0m[38;2;199;183;153m@[0m[38;2;105;88;61mS[0m[38;2;169;152;120m@[0m[38;2;159;143;110m&[0m[38;2;187;172;134m@[0m[38;2;216;201;165m@[0m[38;2;176;159;127m@[0m[38;2;154;134;103m&[0m[38;2;150;127;97m&[0m[38;2;99;77;50mG[0m[38;2;101;82;54mG[0m[38;2;179;163;128m@[0m[38;2;193;181;140m@[0m[38;2;222;207;171m@[0m[38;2;176;160;128m@[0m[38;2;144;127;97mB[0m[38;2;190;174;141m@[0m[38;2;205;189;154m@[0m[38;2;208;192;158m@[0m[38;2;193;177;141m@[0m[38;2;185;170;132m@[0m[38;2;192;177;138m@[0m[38;2;197;181;141m@[0m[38;2;200;186;146m@[0m[38;2;149;135;103m&[0m[38;2;88;71;50mH[0m[38;2;60;38;26m2[0m[38;2;46;19;12ms[0m[38;2;59;13;11ms[0m[38;2;77;8;11mX[0m[38;2;84;7;9mA[0m[38;2;85;8;6mX[0m[38;2;82;8;5mX[0m[38;2;74;7;5mX[0m[38;2;73;14;7mX[0m[38;2;127;78;49mS[0m[38;2;151;108;62m9[0m[38;2;151;110;61m9[0m[38;2;151;109;61m9[0m[38;2;150;108;60m9[0m[38;2;151;109;61m9[0m[38;2;169;127;79m&[0m[38;2;172;131;83m&[0m[38;2;173;133;84m&[0m[38;2;171;132;83m&[0m[38;2;172;134;86m&[0m[38;2;147;111;67m9[0m[38;2;112;78;39mG[0m[38;2;128;91;53m#[0m[38;2;154;112;70mB[0m[38;2;172;130;82m&[0m[38;2;183;145;92m&[0m[38;2;184;149;93m&[0m[38;2;183;149;93m&[0m[38;2;184;148;95m&[0m[38;2;183;149;94m&[0m[38;2;181;148;94m&[0m[38;2;182;148;94m&[0m[38;2;184;148;94m&[0m[38;2;185;147;95m&[0m[38;2;185;148;95m@[0m[38;2;186;149;96m@[0m[38;2;179;141;93m&[0m[38;2;144;106;63m9[0m[38;2;118;79;44mG[0m[38;2;113;74;42mG[0m[38;2;115;75;45mG[0m[38;2;118;78;49mS[0m[38;2;119;79;50mS[0m[38;2;124;81;52mS[0m[38;2;131;87;57m#[0m[38;2;137;90;61m#[0m[38;2;140;92;63m#[0m[38;2;128;82;53mS[0m[38;2;119;77;46mG[0m[38;2;101;64;35mM[0m[38;2;95;63;40mM[0m[38;2;71;44;27m5[0m[38;2;44;26;14ms[0m");
	$display("[38;2;161;122;72mB[0m[38;2;163;123;73mB[0m[38;2;163;123;74mB[0m[38;2;163;124;74mB[0m[38;2;166;126;76mB[0m[38;2;169;128;78m&[0m[38;2;172;131;80m&[0m[38;2;174;133;80m&[0m[38;2;175;134;78m&[0m[38;2;173;134;78m&[0m[38;2;171;134;78m&[0m[38;2;172;134;79m&[0m[38;2;172;135;79m&[0m[38;2;171;135;79m&[0m[38;2;173;134;80m&[0m[38;2;174;134;79m&[0m[38;2;173;134;79m&[0m[38;2;173;134;79m&[0m[38;2;173;133;78m&[0m[38;2;173;134;78m&[0m[38;2;174;134;78m&[0m[38;2;174;135;79m&[0m[38;2;174;135;79m&[0m[38;2;174;135;80m&[0m[38;2;175;135;80m&[0m[38;2;174;135;80m&[0m[38;2;174;135;80m&[0m[38;2;174;135;80m&[0m[38;2;174;135;80m&[0m[38;2;174;135;79m&[0m[38;2;175;135;80m&[0m[38;2;175;136;80m&[0m[38;2;175;136;80m&[0m[38;2;174;135;79m&[0m[38;2;174;135;79m&[0m[38;2;173;134;78m&[0m[38;2;173;134;78m&[0m[38;2;174;133;78m&[0m[38;2;174;133;79m&[0m[38;2;174;133;79m&[0m[38;2;174;133;78m&[0m[38;2;173;133;78m&[0m[38;2;172;134;76m&[0m[38;2;175;128;82m&[0m[38;2;104;48;30mM[0m[38;2;69;19;11mX[0m[38;2;174;142;114m@[0m[38;2;188;165;132m@[0m[38;2;123;106;73m9[0m[38;2;187;169;135m@[0m[38;2;175;155;120m@[0m[38;2;162;147;110m&[0m[38;2;192;176;139m@[0m[38;2;178;163;124m@[0m[38;2;164;149;110m&[0m[38;2;206;190;153m@[0m[38;2;104;87;58mS[0m[38;2;124;106;81m9[0m[38;2;159;142;111m&[0m[38;2;162;145;109m&[0m[38;2;191;174;135m@[0m[38;2;209;194;161m@[0m[38;2;113;97;70m#[0m[38;2;136;116;86mB[0m[38;2;167;139;104m&[0m[38;2;193;161;122m@[0m[38;2;129;101;72m9[0m[38;2;103;81;59mG[0m[38;2;176;163;127m@[0m[38;2;202;187;149m@[0m[38;2;223;207;173m@[0m[38;2;132;115;84m9[0m[38;2;146;130;99m&[0m[38;2;190;175;140m@[0m[38;2;205;190;149m@[0m[38;2;197;182;142m@[0m[38;2;186;171;133m@[0m[38;2;177;161;125m@[0m[38;2;190;174;137m@[0m[38;2;192;176;134m@[0m[38;2;205;186;144m@[0m[38;2;161;142;108m&[0m[38;2;121;102;77m9[0m[38;2;102;87;64mS[0m[38;2;58;41;24m2[0m[38;2;46;16;9mr[0m[38;2;66;10;12mX[0m[38;2;80;7;8mX[0m[38;2;78;7;6mX[0m[38;2;76;5;9mX[0m[38;2;70;3;8ms[0m[38;2;83;25;16m2[0m[38;2;140;96;56m#[0m[38;2;148;108;58m9[0m[38;2;147;107;58m9[0m[38;2;146;106;57m9[0m[38;2;147;107;58m9[0m[38;2;165;125;76mB[0m[38;2;171;131;82m&[0m[38;2;171;132;83m&[0m[38;2;170;132;83m&[0m[38;2;171;133;85m&[0m[38;2;146;112;67m9[0m[38;2;110;78;40mG[0m[38;2;126;90;52mS[0m[38;2;151;110;68m9[0m[38;2;170;127;82m&[0m[38;2;182;142;93m&[0m[38;2;183;147;94m&[0m[38;2;183;146;95m&[0m[38;2;183;146;95m&[0m[38;2;183;147;94m&[0m[38;2;183;147;93m&[0m[38;2;183;147;93m&[0m[38;2;184;145;93m&[0m[38;2;186;146;95m&[0m[38;2;182;142;93m&[0m[38;2;163;122;79mB[0m[38;2;144;102;65m9[0m[38;2;134;91;57m#[0m[38;2;129;85;54mS[0m[38;2;130;86;54m#[0m[38;2;124;80;48mS[0m[38;2;125;80;50mS[0m[38;2;125;81;51mS[0m[38;2;126;81;52mS[0m[38;2;131;87;58m#[0m[38;2;136;93;61m#[0m[38;2;139;97;61m#[0m[38;2;146;103;67m9[0m[38;2;162;119;78mB[0m[38;2;178;136;89m&[0m[38;2;182;141;93m&[0m[38;2;172;131;87m&[0m[38;2;138;100;65m9[0m");
	$display("[38;2;106;76;49mG[0m[38;2;110;78;53mG[0m[38;2;112;78;52mG[0m[38;2;114;81;51mS[0m[38;2;115;83;52mS[0m[38;2;116;82;54mS[0m[38;2;120;86;56mS[0m[38;2;129;93;59m#[0m[38;2;137;101;62m9[0m[38;2;150;114;70mB[0m[38;2;163;125;76mB[0m[38;2;169;131;75m&[0m[38;2;169;132;75m&[0m[38;2;168;132;77m&[0m[38;2;169;131;81m&[0m[38;2;171;132;78m&[0m[38;2;171;132;76m&[0m[38;2;172;131;77m&[0m[38;2;172;132;77m&[0m[38;2;172;133;78m&[0m[38;2;172;133;78m&[0m[38;2;172;133;77m&[0m[38;2;172;133;77m&[0m[38;2;172;133;78m&[0m[38;2;173;134;79m&[0m[38;2;173;134;79m&[0m[38;2;172;133;78m&[0m[38;2;172;133;78m&[0m[38;2;172;133;78m&[0m[38;2;173;134;79m&[0m[38;2;172;133;78m&[0m[38;2;172;133;78m&[0m[38;2;172;133;78m&[0m[38;2;173;134;79m&[0m[38;2;173;134;79m&[0m[38;2;172;133;78m&[0m[38;2;171;132;77m&[0m[38;2;172;131;77m&[0m[38;2;172;131;77m&[0m[38;2;172;131;77m&[0m[38;2;172;131;77m&[0m[38;2;170;130;78m&[0m[38;2;170;130;71mB[0m[38;2;173;129;75m&[0m[38;2;125;83;53mS[0m[38;2;144;111;84mB[0m[38;2;193;173;141m@[0m[38;2;106;89;59mS[0m[38;2;155;140;110m&[0m[38;2;172;155;124m@[0m[38;2;123;105;72m9[0m[38;2;175;158;120m@[0m[38;2;185;168;132m@[0m[38;2;137;120;86mB[0m[38;2;178;160;128m@[0m[38;2;132;114;84m9[0m[38;2;70;51;25m5[0m[38;2;163;145;119m&[0m[38;2;126;109;77m9[0m[38;2;178;162;123m@[0m[38;2;188;173;132m@[0m[38;2;182;165;131m@[0m[38;2;74;59;34mh[0m[38;2;129;111;83m9[0m[38;2;161;132;96m&[0m[38;2;196;161;120m@[0m[38;2;202;172;130m@[0m[38;2;132;108;73m9[0m[38;2;104;87;61mS[0m[38;2;179;164;131m@[0m[38;2;212;197;156m@[0m[38;2;193;177;142m@[0m[38;2;96;79;50mG[0m[38;2;168;152;118m@[0m[38;2;189;174;133m@[0m[38;2;191;176;136m@[0m[38;2;190;175;137m@[0m[38;2;161;145;110m&[0m[38;2;177;162;127m@[0m[38;2;179;164;128m@[0m[38;2;187;171;132m@[0m[38;2;200;184;149m@[0m[38;2;133;117;87mB[0m[38;2;129;111;82m9[0m[38;2;156;142;108m&[0m[38;2;106;93;68mS[0m[38;2;56;29;19mA[0m[38;2;54;9;4mr[0m[38;2;66;8;7ms[0m[38;2;72;5;7ms[0m[38;2;76;5;6mX[0m[38;2;73;7;2ms[0m[38;2;114;65;37mH[0m[38;2;147;106;60m9[0m[38;2;146;105;56m9[0m[38;2;146;104;58m9[0m[38;2;146;105;56m9[0m[38;2;162;124;74mB[0m[38;2;169;131;82m&[0m[38;2;169;131;82m&[0m[38;2;169;131;82m&[0m[38;2;170;132;83m&[0m[38;2;144;109;66m9[0m[38;2;106;76;42mG[0m[38;2;125;87;54mS[0m[38;2;152;110;68m9[0m[38;2;170;126;82m&[0m[38;2;181;139;93m&[0m[38;2;182;144;95m&[0m[38;2;183;145;96m&[0m[38;2;183;144;96m&[0m[38;2;182;144;95m&[0m[38;2;182;145;92m&[0m[38;2;183;146;92m&[0m[38;2;182;145;94m&[0m[38;2;171;132;88m&[0m[38;2;147;105;66m9[0m[38;2;139;97;58m#[0m[38;2;147;104;68m9[0m[38;2;150;106;71m9[0m[38;2;148;102;66m9[0m[38;2;148;102;69m9[0m[38;2;144;99;67m9[0m[38;2;142;97;65m9[0m[38;2;139;95;63m#[0m[38;2;144;99;66m9[0m[38;2;159;115;78mB[0m[38;2;172;131;89m&[0m[38;2;182;142;95m&[0m[38;2;185;145;96m&[0m[38;2;185;144;96m&[0m[38;2;184;143;94m&[0m[38;2;183;143;94m&[0m[38;2;183;142;93m&[0m[38;2;177;136;87m&[0m");
	$display("[38;2;105;75;49mG[0m[38;2;111;77;53mG[0m[38;2;119;83;60mS[0m[38;2;122;87;60mS[0m[38;2;121;87;59mS[0m[38;2;117;84;58mS[0m[38;2;114;81;56mS[0m[38;2;111;78;53mG[0m[38;2;108;76;47mG[0m[38;2;111;77;48mG[0m[38;2;125;90;55m#[0m[38;2;142;104;62m9[0m[38;2;158;121;74mB[0m[38;2;166;129;81m&[0m[38;2;167;130;78m&[0m[38;2;169;129;75m&[0m[38;2;169;130;74m&[0m[38;2;170;129;75m&[0m[38;2;169;129;77m&[0m[38;2;169;129;77m&[0m[38;2;169;129;77m&[0m[38;2;169;129;78m&[0m[38;2;169;129;78m&[0m[38;2;169;130;77m&[0m[38;2;170;130;77m&[0m[38;2;170;130;77m&[0m[38;2;170;130;77m&[0m[38;2;170;130;77m&[0m[38;2;170;130;77m&[0m[38;2;171;131;78m&[0m[38;2;170;131;78m&[0m[38;2;169;130;77m&[0m[38;2;169;130;77m&[0m[38;2;169;130;77m&[0m[38;2;169;129;76m&[0m[38;2;169;129;76m&[0m[38;2;168;129;76m&[0m[38;2;170;129;76m&[0m[38;2;170;129;76m&[0m[38;2;170;129;76m&[0m[38;2;170;129;76m&[0m[38;2;170;128;75m&[0m[38;2;168;127;74mB[0m[38;2;164;127;77mB[0m[38;2;155;127;83mB[0m[38;2;183;164;125m@[0m[38;2;125;109;83m9[0m[38;2;100;84;59mG[0m[38;2;171;153;128m@[0m[38;2;107;89;65mS[0m[38;2;108;92;64mS[0m[38;2;183;168;130m@[0m[38;2;155;138;105m&[0m[38;2;117;99;71m#[0m[38;2;154;136;111m&[0m[38;2;54;36;16mA[0m[38;2;108;91;70mS[0m[38;2;132;116;90mB[0m[38;2;124;108;75m9[0m[38;2;183;169;132m@[0m[38;2;182;168;129m@[0m[38;2;150;131;99m&[0m[38;2;82;63;39mM[0m[38;2;136;118;89mB[0m[38;2;156;130;94m&[0m[38;2;194;160;121m@[0m[38;2;204;170;123m@[0m[38;2;201;171;127m@[0m[38;2;127;105;73m9[0m[38;2;111;93;66m#[0m[38;2;184;169;131m@[0m[38;2;210;195;156m@[0m[38;2;123;106;78m9[0m[38;2;103;86;59mS[0m[38;2;184;168;133m@[0m[38;2;186;170;131m@[0m[38;2;186;172;132m@[0m[38;2;174;158;123m@[0m[38;2;145;129;97mB[0m[38;2;172;155;124m@[0m[38;2;148;132;98m&[0m[38;2;188;172;135m@[0m[38;2;192;177;139m@[0m[38;2;102;84;56mG[0m[38;2;136;113;84mB[0m[38;2;184;166;126m@[0m[38;2;158;145;109m&[0m[38;2;83;64;43mM[0m[38;2;52;15;8ms[0m[38;2;65;8;7ms[0m[38;2;76;6;8mX[0m[38;2;76;5;5mX[0m[38;2;91;40;22m3[0m[38;2;141;100;61m9[0m[38;2;142;103;53m#[0m[38;2;143;103;56m9[0m[38;2;143;104;55m9[0m[38;2;160;122;73mB[0m[38;2;168;130;81m&[0m[38;2;168;130;81m&[0m[38;2;168;130;81m&[0m[38;2;169;130;81m&[0m[38;2;143;108;65m9[0m[38;2;105;75;41mH[0m[38;2;124;86;53mS[0m[38;2;150;108;66m9[0m[38;2;167;124;79mB[0m[38;2;178;139;92m&[0m[38;2;180;144;95m&[0m[38;2;181;145;95m&[0m[38;2;180;143;93m&[0m[38;2;180;142;91m&[0m[38;2;180;143;90m&[0m[38;2;180;143;93m&[0m[38;2;161;123;80mB[0m[38;2;140;99;62m9[0m[38;2;146;102;68m9[0m[38;2;158;114;77mB[0m[38;2;164;119;81mB[0m[38;2;158;113;74mB[0m[38;2;149;104;66m9[0m[38;2;149;104;68m9[0m[38;2;147;103;69m9[0m[38;2;148;104;68m9[0m[38;2;157;114;76mB[0m[38;2;174;130;92m&[0m[38;2;185;142;101m@[0m[38;2;186;145;99m@[0m[38;2;186;145;96m&[0m[38;2;184;146;95m&[0m[38;2;182;143;94m&[0m[38;2;182;143;94m&[0m[38;2;181;142;93m&[0m[38;2;179;140;92m&[0m[38;2;172;131;85m&[0m");
	$display("[38;2;158;117;86mB[0m[38;2;144;104;74m9[0m[38;2;129;92;64m#[0m[38;2;119;83;57mS[0m[38;2;116;83;57mS[0m[38;2;117;85;58mS[0m[38;2;119;85;58mS[0m[38;2;125;91;61m#[0m[38;2;126;91;58m#[0m[38;2;125;90;56m#[0m[38;2;122;86;57mS[0m[38;2;121;84;57mS[0m[38;2;125;88;56mS[0m[38;2;140;104;64m9[0m[38;2;160;124;75mB[0m[38;2;168;129;73mB[0m[38;2;168;127;74mB[0m[38;2;168;127;76mB[0m[38;2;167;127;75mB[0m[38;2;168;126;76mB[0m[38;2;167;126;76mB[0m[38;2;167;126;76mB[0m[38;2;167;126;76mB[0m[38;2;166;127;75mB[0m[38;2;166;127;75mB[0m[38;2;166;127;75mB[0m[38;2;167;128;76mB[0m[38;2;168;128;76m&[0m[38;2;168;128;76m&[0m[38;2;168;128;76m&[0m[38;2;168;128;75mB[0m[38;2;167;128;74mB[0m[38;2;167;127;75mB[0m[38;2;167;127;75mB[0m[38;2;167;126;75mB[0m[38;2;167;127;75mB[0m[38;2;168;127;75mB[0m[38;2;168;127;75mB[0m[38;2;167;126;74mB[0m[38;2;167;126;74mB[0m[38;2;167;126;74mB[0m[38;2;168;125;74mB[0m[38;2;168;126;76mB[0m[38;2;155;122;77mB[0m[38;2;169;145;105m&[0m[38;2;166;146;115m&[0m[38;2;71;54;33m3[0m[38;2;132;116;91mB[0m[38;2;117;100;80m#[0m[38;2;50;35;16mA[0m[38;2;137;124;95mB[0m[38;2;178;163;129m@[0m[38;2;103;89;61mS[0m[38;2;129;117;88mB[0m[38;2;75;61;42mh[0m[38;2;53;37;22mA[0m[38;2;127;112;88m9[0m[38;2;73;58;33mh[0m[38;2;140;125;99mB[0m[38;2;181;166;129m@[0m[38;2;176;161;123m@[0m[38;2;114;91;64mS[0m[38;2;121;96;71m#[0m[38;2;148;124;93mB[0m[38;2;149;123;89mB[0m[38;2;195;163;124m@[0m[38;2;203;168;123m@[0m[38;2;202;170;126m@[0m[38;2;194;169;125m@[0m[38;2;120;99;62m#[0m[38;2;120;100;72m#[0m[38;2;190;174;139m@[0m[38;2;167;151;117m@[0m[38;2;70;52;33m3[0m[38;2;152;136;107m&[0m[38;2;185;169;132m@[0m[38;2;183;168;127m@[0m[38;2;186;170;134m@[0m[38;2;132;115;84m9[0m[38;2;170;154;123m@[0m[38;2;131;114;83m9[0m[38;2;149;133;99m&[0m[38;2;192;177;136m@[0m[38;2;164;148;116m@[0m[38;2;79;60;38mh[0m[38;2;146;132;98m&[0m[38;2;186;173;129m@[0m[38;2;181;166;128m@[0m[38;2;104;84;60mS[0m[38;2;59;18;13mX[0m[38;2;73;8;9mX[0m[38;2;74;6;8mX[0m[38;2;78;28;18m2[0m[38;2;136;94;59m#[0m[38;2;140;101;53m#[0m[38;2;140;102;54m#[0m[38;2;140;102;54m#[0m[38;2;159;121;73mB[0m[38;2;167;129;81m&[0m[38;2;166;128;80m&[0m[38;2;167;129;81m&[0m[38;2;167;129;81m&[0m[38;2;141;109;63m9[0m[38;2;102;74;39mH[0m[38;2;120;84;50mS[0m[38;2;146;107;65m9[0m[38;2;165;124;78mB[0m[38;2;176;138;91m&[0m[38;2;179;143;94m&[0m[38;2;179;143;93m&[0m[38;2;179;143;92m&[0m[38;2;180;144;92m&[0m[38;2;177;140;92m&[0m[38;2;153;114;71mB[0m[38;2;138;99;59m#[0m[38;2;152;110;71mB[0m[38;2;162;118;79mB[0m[38;2;164;119;80mB[0m[38;2;164;119;80mB[0m[38;2;156;112;72mB[0m[38;2;148;102;63m9[0m[38;2;147;102;64m9[0m[38;2;154;110;70mB[0m[38;2;169;126;85m&[0m[38;2;182;139;97m&[0m[38;2;184;141;98m&[0m[38;2;183;141;96m&[0m[38;2;182;142;97m&[0m[38;2;183;143;99m&[0m[38;2;183;143;100m&[0m[38;2;183;142;98m&[0m[38;2;182;142;96m&[0m[38;2;182;141;95m&[0m[38;2;180;139;93m&[0m[38;2;181;140;93m&[0m");
	$display("[38;2;167;125;94m&[0m[38;2;169;128;95m&[0m[38;2;167;129;95m&[0m[38;2;158;121;90mB[0m[38;2;138;103;74m9[0m[38;2;124;90;60m#[0m[38;2;129;93;62m#[0m[38;2;145;106;74m9[0m[38;2;148;106;73m9[0m[38;2;147;106;70m9[0m[38;2;141;101;67m9[0m[38;2;131;93;62m#[0m[38;2;122;86;56mS[0m[38;2;120;85;52mS[0m[38;2;127;91;56m#[0m[38;2;151;113;71mB[0m[38;2;163;125;77mB[0m[38;2;163;125;73mB[0m[38;2;165;124;74mB[0m[38;2;165;124;76mB[0m[38;2;165;124;75mB[0m[38;2;164;125;74mB[0m[38;2;164;125;74mB[0m[38;2;165;125;74mB[0m[38;2;165;125;74mB[0m[38;2;166;125;75mB[0m[38;2;166;126;77mB[0m[38;2;167;126;77mB[0m[38;2;166;126;74mB[0m[38;2;166;125;74mB[0m[38;2;165;125;74mB[0m[38;2;165;125;72mB[0m[38;2;165;125;72mB[0m[38;2;165;125;72mB[0m[38;2;165;125;72mB[0m[38;2;165;125;72mB[0m[38;2;164;125;72mB[0m[38;2;164;125;72mB[0m[38;2;164;124;71mB[0m[38;2;164;124;71mB[0m[38;2;164;124;71mB[0m[38;2;164;124;72mB[0m[38;2;161;124;74mB[0m[38;2;151;125;79mB[0m[38;2;177;159;123m@[0m[38;2;114;99;73m#[0m[38;2;62;52;35m3[0m[38;2;105;94;74m#[0m[38;2;50;35;23mA[0m[38;2;60;43;28m5[0m[38;2;161;144;112m&[0m[38;2;151;132;104m&[0m[38;2;85;68;51mH[0m[38;2;97;82;61mG[0m[38;2;45;28;17mX[0m[38;2;79;62;52mM[0m[38;2;82;67;50mM[0m[38;2;56;41;23m2[0m[38;2;134;118;91mB[0m[38;2;183;166;130m@[0m[38;2;149;134;100m&[0m[38;2;100;79;53mG[0m[38;2;156;130;101m&[0m[38;2;142;118;88mB[0m[38;2;141;117;86mB[0m[38;2;194;164;124m@[0m[38;2;199;167;121m@[0m[38;2;202;168;124m@[0m[38;2;203;170;121m@[0m[38;2;196;167;119m@[0m[38;2;116;90;58mS[0m[38;2;131;112;80m9[0m[38;2;179;164;130m@[0m[38;2;88;72;50mH[0m[38;2;103;88;62mS[0m[38;2;182;166;132m@[0m[38;2;181;167;127m@[0m[38;2;185;169;133m@[0m[38;2;142;125;92mB[0m[38;2;144;128;93mB[0m[38;2;168;152;120m@[0m[38;2;98;81;52mG[0m[38;2;170;154;117m@[0m[38;2;191;175;136m@[0m[38;2;104;88;63mS[0m[38;2;93;76;55mG[0m[38;2;173;158;123m@[0m[38;2;189;173;128m@[0m[38;2;175;161;122m@[0m[38;2;93;71;49mH[0m[38;2;64;12;9ms[0m[38;2;72;4;9ms[0m[38;2;84;34;22m5[0m[38;2;135;95;60m#[0m[38;2;136;98;53m#[0m[38;2;137;98;55m#[0m[38;2;137;99;54m#[0m[38;2;156;118;72mB[0m[38;2;166;128;81m&[0m[38;2;165;127;81m&[0m[38;2;166;128;82m&[0m[38;2;166;129;81m&[0m[38;2;141;109;65m9[0m[38;2;100;72;38mH[0m[38;2;117;81;49mS[0m[38;2;143;104;64m9[0m[38;2;162;121;76mB[0m[38;2;175;137;89m&[0m[38;2;177;141;90m&[0m[38;2;178;141;91m&[0m[38;2;178;142;92m&[0m[38;2;174;139;91m&[0m[38;2;146;109;66m9[0m[38;2;140;102;62m9[0m[38;2;154;115;76mB[0m[38;2;160;120;80mB[0m[38;2;161;117;78mB[0m[38;2;162;117;78mB[0m[38;2;163;118;79mB[0m[38;2;156;112;73mB[0m[38;2;151;107;67m9[0m[38;2;169;124;84m&[0m[38;2;180;137;95m&[0m[38;2;182;140;97m&[0m[38;2;182;140;96m&[0m[38;2;181;140;94m&[0m[38;2;180;139;94m&[0m[38;2;181;139;95m&[0m[38;2;181;139;96m&[0m[38;2;181;138;96m&[0m[38;2;182;139;95m&[0m[38;2;181;140;94m&[0m[38;2;182;140;95m&[0m[38;2;178;136;95m&[0m[38;2;163;120;87mB[0m");
	$display("[38;2;165;124;93m&[0m[38;2;168;127;93m&[0m[38;2;170;130;95m&[0m[38;2;170;131;95m&[0m[38;2;170;130;95m&[0m[38;2;165;124;90m&[0m[38;2;157;116;82mB[0m[38;2;148;108;73m9[0m[38;2;146;105;70m9[0m[38;2;147;107;71m9[0m[38;2;147;106;70m9[0m[38;2;146;107;71m9[0m[38;2;141;103;68m9[0m[38;2;131;93;59m#[0m[38;2;121;84;55mS[0m[38;2;118;82;54mS[0m[38;2;135;101;60m#[0m[38;2;159;122;76mB[0m[38;2;173;132;88m&[0m[38;2;178;137;91m&[0m[38;2;177;137;89m&[0m[38;2;175;138;87m&[0m[38;2;174;138;85m&[0m[38;2;173;136;85m&[0m[38;2;171;134;85m&[0m[38;2;167;130;84m&[0m[38;2;150;113;70mB[0m[38;2;150;112;67m9[0m[38;2;161;122;73mB[0m[38;2;162;123;73mB[0m[38;2;163;124;73mB[0m[38;2;162;123;72mB[0m[38;2;162;123;73mB[0m[38;2;161;122;73mB[0m[38;2;160;122;72mB[0m[38;2;161;122;72mB[0m[38;2;161;123;73mB[0m[38;2;161;122;73mB[0m[38;2;160;121;71mB[0m[38;2;160;121;72mB[0m[38;2;160;121;72mB[0m[38;2;160;121;72mB[0m[38;2;155;120;72mB[0m[38;2;157;133;90m&[0m[38;2;168;151;120m@[0m[38;2;68;54;35m3[0m[38;2;55;41;31m2[0m[38;2;47;34;21mA[0m[38;2;54;35;26m2[0m[38;2;107;87;70mS[0m[38;2;159;143;110m&[0m[38;2;89;72;55mH[0m[38;2;68;51;43m3[0m[38;2;50;35;22mA[0m[38;2;48;33;22mA[0m[38;2;65;50;40m3[0m[38;2;44;31;22mX[0m[38;2;50;36;22mA[0m[38;2;141;125;94mB[0m[38;2;178;160;127m@[0m[38;2;98;80;53mG[0m[38;2;131;106;77m9[0m[38;2;167;139;109m&[0m[38;2;130;102;76m9[0m[38;2;134;106;79m9[0m[38;2;179;151;113m@[0m[38;2;174;146;106m&[0m[38;2;173;142;104m&[0m[38;2;176;145;104m&[0m[38;2;181;150;107m@[0m[38;2;175;147;112m@[0m[38;2;99;76;49mG[0m[38;2;148;130;103m&[0m[38;2;121;104;78m9[0m[38;2;68;52;31m3[0m[38;2;169;153;121m@[0m[38;2;182;166;127m@[0m[38;2;183;166;129m@[0m[38;2;151;133;105m&[0m[38;2;106;89;63mS[0m[38;2;182;165;132m@[0m[38;2;117;99;74m#[0m[38;2;108;92;64mS[0m[38;2;182;167;130m@[0m[38;2;152;137;103m&[0m[38;2;64;48;27m5[0m[38;2;144;128;104m&[0m[38;2;184;167;128m@[0m[38;2;187;172;129m@[0m[38;2;166;145;112m&[0m[38;2;75;32;25m5[0m[38;2;57;4;3mr[0m[38;2;103;62;37mH[0m[38;2;134;98;57m#[0m[38;2;134;97;53m#[0m[38;2;135;97;54m#[0m[38;2;137;98;54m#[0m[38;2;155;116;72mB[0m[38;2;165;127;82m&[0m[38;2;165;126;81m&[0m[38;2;165;126;82m&[0m[38;2;166;128;81m&[0m[38;2;141;109;66m9[0m[38;2;99;72;39mH[0m[38;2;115;79;49mG[0m[38;2;141;101;63m9[0m[38;2;159;118;76mB[0m[38;2;173;135;85m&[0m[38;2;175;140;85m&[0m[38;2;177;142;92m&[0m[38;2;171;134;88m&[0m[38;2;144;104;62m9[0m[38;2;144;103;65m9[0m[38;2;160;117;82mB[0m[38;2;162;119;83mB[0m[38;2;160;117;79mB[0m[38;2;160;117;78mB[0m[38;2;160;115;77mB[0m[38;2;161;117;78mB[0m[38;2;168;124;85m&[0m[38;2;178;136;94m&[0m[38;2;182;140;97m&[0m[38;2;180;139;95m&[0m[38;2;180;139;94m&[0m[38;2;179;139;95m&[0m[38;2;178;139;95m&[0m[38;2;179;138;95m&[0m[38;2;179;139;93m&[0m[38;2;180;139;90m&[0m[38;2;181;137;90m&[0m[38;2;181;138;92m&[0m[38;2;176;135;93m&[0m[38;2;157;117;84mB[0m[38;2;122;83;57mS[0m[38;2;105;68;45mH[0m");
	$display("[38;2;163;123;88m&[0m[38;2;164;124;89m&[0m[38;2;166;125;90m&[0m[38;2;166;126;91m&[0m[38;2;166;126;91m&[0m[38;2;168;128;92m&[0m[38;2;168;128;93m&[0m[38;2;165;125;90m&[0m[38;2;157;117;82mB[0m[38;2;147;107;72m9[0m[38;2;144;104;69m9[0m[38;2;145;105;70m9[0m[38;2;145;105;70m9[0m[38;2;145;105;70m9[0m[38;2;139;100;65m9[0m[38;2;127;91;59m#[0m[38;2;117;82;50mS[0m[38;2;129;91;56m#[0m[38;2;173;132;93m&[0m[38;2;191;152;102m@[0m[38;2;186;148;96m@[0m[38;2;183;145;97m&[0m[38;2;181;144;95m&[0m[38;2;180;143;94m&[0m[38;2;168;131;86m&[0m[38;2;149;113;74mB[0m[38;2;135;101;64m9[0m[38;2;119;84;45mS[0m[38;2;151;113;68mB[0m[38;2;157;119;71mB[0m[38;2;157;120;69mB[0m[38;2;158;120;71mB[0m[38;2;157;120;71mB[0m[38;2;157;119;70mB[0m[38;2;158;120;71mB[0m[38;2;158;120;71mB[0m[38;2;157;119;70mB[0m[38;2;157;119;69mB[0m[38;2;157;119;69mB[0m[38;2;157;119;69mB[0m[38;2;157;119;69mB[0m[38;2;157;120;69mB[0m[38;2;149;116;67mB[0m[38;2;165;141;98m&[0m[38;2;143;126;98mB[0m[38;2;45;30;18mX[0m[38;2;40;26;19ms[0m[38;2;42;28;16mX[0m[38;2;98;75;59mG[0m[38;2;134;113;89mB[0m[38;2;123;112;86m9[0m[38;2;45;31;18mX[0m[38;2;45;28;22mX[0m[38;2;46;29;21mX[0m[38;2;45;29;21mX[0m[38;2;45;29;23mX[0m[38;2;41;28;20mX[0m[38;2;65;52;32m3[0m[38;2;169;149;121m@[0m[38;2;127;106;83m9[0m[38;2;76;54;34mh[0m[38;2;183;152;110m@[0m[38;2;168;141;103m&[0m[38;2;108;83;59mS[0m[38;2;153;121;90mB[0m[38;2;199;166;124m@[0m[38;2;196;164;119m@[0m[38;2;193;161;116m@[0m[38;2;190;158;114m@[0m[38;2;185;153;107m@[0m[38;2;178;148;106m@[0m[38;2;152;124;90mB[0m[38;2;96;75;50mH[0m[38;2;122;106;88m9[0m[38;2;54;38;24m2[0m[38;2;143;126;98mB[0m[38;2;182;164;126m@[0m[38;2;181;164;125m@[0m[38;2;154;138;105m&[0m[38;2;58;42;27m2[0m[38;2;134;117;90mB[0m[38;2;165;145;115m&[0m[38;2;69;54;35m3[0m[38;2;145;132;101m&[0m[38;2;172;156;123m@[0m[38;2;73;59;38mh[0m[38;2;98;84;62mG[0m[38;2;178;162;124m@[0m[38;2;184;170;123m@[0m[38;2;183;167;126m@[0m[38;2;130;103;79m9[0m[38;2;78;40;23m5[0m[38;2;128;92;56m#[0m[38;2;131;98;54m#[0m[38;2;131;97;52m#[0m[38;2;133;96;52m#[0m[38;2;134;95;53m#[0m[38;2;153;113;70mB[0m[38;2;163;124;80mB[0m[38;2;163;124;80mB[0m[38;2;163;124;79mB[0m[38;2;163;125;78mB[0m[38;2;140;109;67m9[0m[38;2;97;71;38mH[0m[38;2;111;77;46mG[0m[38;2;139;100;61m9[0m[38;2;156;117;74mB[0m[38;2;169;133;81m&[0m[38;2;173;137;87m&[0m[38;2;166;128;88m&[0m[38;2;137;100;62m9[0m[38;2;144;103;68m9[0m[38;2;159;115;80mB[0m[38;2;160;116;79mB[0m[38;2;160;116;78mB[0m[38;2;159;116;79mB[0m[38;2;159;115;79mB[0m[38;2;165;121;83mB[0m[38;2;176;132;92m&[0m[38;2;182;138;97m&[0m[38;2;180;138;95m&[0m[38;2;180;138;96m&[0m[38;2;179;138;95m&[0m[38;2;179;138;94m&[0m[38;2;179;138;94m&[0m[38;2;179;138;94m&[0m[38;2;178;139;91m&[0m[38;2;179;139;91m&[0m[38;2;181;138;91m&[0m[38;2;172;130;88m&[0m[38;2;147;108;72m9[0m[38;2;114;78;50mG[0m[38;2;101;65;42mH[0m[38;2;110;73;49mG[0m[38;2;125;84;54mS[0m");
	$display("[38;2;161;121;86mB[0m[38;2;162;121;86mB[0m[38;2;163;123;88m&[0m[38;2;163;123;88m&[0m[38;2;164;124;89m&[0m[38;2;165;125;90m&[0m[38;2;165;125;90m&[0m[38;2;166;126;91m&[0m[38;2;167;127;92m&[0m[38;2;164;124;89m&[0m[38;2;154;114;79mB[0m[38;2;144;104;69m9[0m[38;2;142;102;67m9[0m[38;2;144;103;68m9[0m[38;2;145;103;68m9[0m[38;2;143;103;70m9[0m[38;2;135;96;65m#[0m[38;2;121;82;54mS[0m[38;2;131;93;63m#[0m[38;2;169;132;91m&[0m[38;2;183;147;96m&[0m[38;2;185;147;98m@[0m[38;2;183;145;95m&[0m[38;2;183;145;96m&[0m[38;2;164;127;82m&[0m[38;2;141;107;67m9[0m[38;2;131;100;62m#[0m[38;2;113;81;41mG[0m[38;2;148;109;64m9[0m[38;2;156;118;70mB[0m[38;2;156;118;67mB[0m[38;2;155;117;68mB[0m[38;2;155;117;68mB[0m[38;2;155;117;68mB[0m[38;2;155;117;68mB[0m[38;2;155;117;68mB[0m[38;2;154;116;67mB[0m[38;2;154;116;68mB[0m[38;2;154;116;68mB[0m[38;2;154;116;68mB[0m[38;2;154;116;68mB[0m[38;2;154;117;70mB[0m[38;2;146;114;70m9[0m[38;2;170;149;110m@[0m[38;2;114;101;76m#[0m[38;2;34;25;15ms[0m[38;2;38;24;17ms[0m[38;2;101;73;55mG[0m[38;2;160;131;99m&[0m[38;2;141;120;92mB[0m[38;2;74;57;39mh[0m[38;2;39;24;13ms[0m[38;2;46;26;21mX[0m[38;2;63;40;31m5[0m[38;2;82;59;48mM[0m[38;2;63;42;31m5[0m[38;2;46;32;18mX[0m[38;2;94;79;60mG[0m[38;2;134;112;91mB[0m[38;2;56;34;20mA[0m[38;2;125;101;79m9[0m[38;2;199;165;124m@[0m[38;2;160;129;96m&[0m[38;2;97;68;47mH[0m[38;2;173;139;108m&[0m[38;2;198;164;120m@[0m[38;2;197;164;118m@[0m[38;2;197;164;117m@[0m[38;2;198;164;119m@[0m[38;2;198;165;118m@[0m[38;2;199;165;116m@[0m[38;2;200;165;122m@[0m[38;2;152;123;93mB[0m[38;2;85;64;47mM[0m[38;2;50;36;23mA[0m[38;2;113;97;73m#[0m[38;2;177;161;127m@[0m[38;2;178;163;123m@[0m[38;2;154;139;104m&[0m[38;2;88;76;52mH[0m[38;2;59;46;33m5[0m[38;2;151;136;107m&[0m[38;2;102;89;65mS[0m[38;2;82;69;46mM[0m[38;2;174;156;126m@[0m[38;2;97;81;57mG[0m[38;2;68;53;32m3[0m[38;2;168;153;119m@[0m[38;2;178;165;119m@[0m[38;2;178;166;121m@[0m[38;2;172;153;115m@[0m[38;2;129;102;64m#[0m[38;2;128;97;52m#[0m[38;2;129;97;51m#[0m[38;2;129;95;53m#[0m[38;2;129;94;52m#[0m[38;2;130;93;50m#[0m[38;2;148;111;67m9[0m[38;2;160;122;77mB[0m[38;2;161;123;78mB[0m[38;2;161;124;78mB[0m[38;2;161;124;77mB[0m[38;2;139;107;66m9[0m[38;2;95;69;38mH[0m[38;2;110;75;47mG[0m[38;2;138;98;61m#[0m[38;2;152;115;74mB[0m[38;2;167;131;86m&[0m[38;2;158;121;80mB[0m[38;2;133;93;60m#[0m[38;2;141;102;67m9[0m[38;2;157;116;80mB[0m[38;2;159;115;80mB[0m[38;2;158;114;77mB[0m[38;2;157;114;76mB[0m[38;2;160;117;80mB[0m[38;2;171;128;89m&[0m[38;2;179;137;97m&[0m[38;2;180;138;96m&[0m[38;2;179;138;94m&[0m[38;2;179;138;94m&[0m[38;2;179;138;95m&[0m[38;2;179;137;95m&[0m[38;2;178;136;94m&[0m[38;2;180;138;94m&[0m[38;2;180;138;94m&[0m[38;2;177;134;93m&[0m[38;2;160;119;84mB[0m[38;2;133;94;65m#[0m[38;2;106;68;44mH[0m[38;2;99;60;38mM[0m[38;2;112;73;50mG[0m[38;2;125;83;55mS[0m[38;2;129;85;52mS[0m[38;2;135;90;55m#[0m");
	$display("[38;2;145;108;80mB[0m[38;2;158;118;87mB[0m[38;2;162;119;86mB[0m[38;2;163;119;85mB[0m[38;2;163;120;86mB[0m[38;2;163;122;88m&[0m[38;2;163;122;90m&[0m[38;2;163;123;89m&[0m[38;2;163;125;88m&[0m[38;2;164;124;89m&[0m[38;2;166;126;91m&[0m[38;2;161;121;86mB[0m[38;2;152;112;77mB[0m[38;2;144;103;69m9[0m[38;2;144;100;67m9[0m[38;2;145;102;70m9[0m[38;2;143;103;72m9[0m[38;2;136;99;69m9[0m[38;2;127;89;63m#[0m[38;2;128;91;60m#[0m[38;2;162;128;84m&[0m[38;2;186;150;99m@[0m[38;2;185;148;95m@[0m[38;2;185;148;96m@[0m[38;2;161;125;80mB[0m[38;2;138;104;65m9[0m[38;2;128;97;58m#[0m[38;2;111;79;40mG[0m[38;2;146;109;64m9[0m[38;2;152;116;65mB[0m[38;2;153;116;68mB[0m[38;2;153;115;66mB[0m[38;2;153;115;66mB[0m[38;2;154;115;66mB[0m[38;2;154;115;67mB[0m[38;2;153;114;66mB[0m[38;2;152;114;66mB[0m[38;2;151;113;68mB[0m[38;2;151;113;68mB[0m[38;2;151;113;68mB[0m[38;2;151;113;68mB[0m[38;2;151;113;67m9[0m[38;2;145;110;74m9[0m[38;2;171;149;114m@[0m[38;2;88;79;55mG[0m[38;2;33;20;14mr[0m[38;2;80;53;41mh[0m[38;2;180;145;107m@[0m[38;2;179;145;101m&[0m[38;2;144;114;89mB[0m[38;2;72;47;31m3[0m[38;2;75;52;38mh[0m[38;2;98;71;50mH[0m[38;2;166;134;106m&[0m[38;2;138;102;74m9[0m[38;2;167;133;101m&[0m[38;2;155;124;90mB[0m[38;2;153;121;89mB[0m[38;2;136;104;74m9[0m[38;2;129;97;68m#[0m[38;2;186;156;114m@[0m[38;2;196;163;122m@[0m[38;2;167;133;99m&[0m[38;2;142;108;75m9[0m[38;2;189;155;117m@[0m[38;2;194;161;119m@[0m[38;2;195;163;119m@[0m[38;2;195;163;119m@[0m[38;2;195;163;119m@[0m[38;2;196;162;118m@[0m[38;2;197;163;118m@[0m[38;2;197;162;116m@[0m[38;2;195;163;122m@[0m[38;2;117;95;66m#[0m[38;2;41;25;10ms[0m[38;2;92;77;60mG[0m[38;2;175;158;121m@[0m[38;2;178;162;121m@[0m[38;2;145;131;101m&[0m[38;2;102;90;67mS[0m[38;2;68;56;43mh[0m[38;2;66;54;35m3[0m[38;2;128;118;93mB[0m[38;2;54;42;25m2[0m[38;2;139;120;98mB[0m[38;2;114;97;73m#[0m[38;2;50;35;21mA[0m[38;2;151;137;107m&[0m[38;2;177;161;122m@[0m[38;2;177;161;120m@[0m[38;2;180;160;120m@[0m[38;2;146;121;84mB[0m[38;2;124;94;52m#[0m[38;2;127;94;51m#[0m[38;2;125;92;51mS[0m[38;2;126;91;51mS[0m[38;2;128;90;51mS[0m[38;2;146;109;67m9[0m[38;2;159;122;78mB[0m[38;2;160;123;78mB[0m[38;2;161;124;79mB[0m[38;2;162;124;79mB[0m[38;2;140;108;65m9[0m[38;2;93;69;34mM[0m[38;2;108;75;45mG[0m[38;2;135;97;61m#[0m[38;2;150;112;75mB[0m[38;2;147;108;71m9[0m[38;2;131;92;56m#[0m[38;2;145;103;69m9[0m[38;2;156;114;78mB[0m[38;2;156;114;78mB[0m[38;2;155;112;76mB[0m[38;2;159;117;80mB[0m[38;2;167;127;89m&[0m[38;2;177;135;97m&[0m[38;2;179;137;97m&[0m[38;2;178;136;95m&[0m[38;2;178;137;93m&[0m[38;2;178;137;92m&[0m[38;2;178;137;93m&[0m[38;2;179;138;93m&[0m[38;2;178;137;93m&[0m[38;2;176;136;94m&[0m[38;2;166;124;87m&[0m[38;2;143;101;71m9[0m[38;2;116;76;52mG[0m[38;2;97;60;39mM[0m[38;2;101;65;44mH[0m[38;2;112;73;51mG[0m[38;2;117;76;50mG[0m[38;2;128;84;54mS[0m[38;2;130;86;55m#[0m[38;2;133;89;59m#[0m[38;2;137;93;60m#[0m");
	$display("[38;2;81;54;38mh[0m[38;2;101;71;55mG[0m[38;2;129;93;74m#[0m[38;2;150;109;84mB[0m[38;2;160;118;87mB[0m[38;2;162;121;86mB[0m[38;2;162;121;86mB[0m[38;2;162;122;87mB[0m[38;2;162;122;87mB[0m[38;2;162;122;87mB[0m[38;2;164;124;89m&[0m[38;2;165;125;90m&[0m[38;2;166;126;91m&[0m[38;2;161;121;86mB[0m[38;2;152;110;75mB[0m[38;2;146;103;70m9[0m[38;2;144;101;69m9[0m[38;2;144;101;70m9[0m[38;2;147;105;75m9[0m[38;2;132;94;63m#[0m[38;2;125;89;55mS[0m[38;2;152;116;76mB[0m[38;2;178;141;95m&[0m[38;2;181;147;95m&[0m[38;2;151;118;74mB[0m[38;2;132;98;63m#[0m[38;2;125;92;60m#[0m[38;2;111;77;43mG[0m[38;2;145;108;65m9[0m[38;2;149;113;65m9[0m[38;2;151;113;68mB[0m[38;2;150;112;66m9[0m[38;2;150;112;66m9[0m[38;2;150;112;67m9[0m[38;2;150;112;67m9[0m[38;2;150;112;67m9[0m[38;2;150;112;67m9[0m[38;2;150;112;67m9[0m[38;2;150;112;67m9[0m[38;2;150;112;67m9[0m[38;2;150;112;67m9[0m[38;2;148;111;65m9[0m[38;2;151;119;79mB[0m[38;2;167;150;111m@[0m[38;2;72;62;44mh[0m[38;2;52;31;21mA[0m[38;2;164;129;100m&[0m[38;2;196;160;113m@[0m[38;2;197;162;109m@[0m[38;2;195;158;115m@[0m[38;2;181;145;107m@[0m[38;2;188;153;114m@[0m[38;2;194;160;116m@[0m[38;2;196;162;115m@[0m[38;2;197;162;115m@[0m[38;2;197;162;116m@[0m[38;2;198;164;117m@[0m[38;2;198;164;115m@[0m[38;2;198;164;118m@[0m[38;2;199;165;120m@[0m[38;2;195;162;116m@[0m[38;2;194;161;116m@[0m[38;2;194;161;117m@[0m[38;2;189;156;112m@[0m[38;2;194;161;116m@[0m[38;2;194;162;116m@[0m[38;2;187;154;112m@[0m[38;2;186;152;111m@[0m[38;2;189;156;113m@[0m[38;2;194;159;118m@[0m[38;2;195;163;121m@[0m[38;2;197;163;114m@[0m[38;2;197;163;115m@[0m[38;2;181;153;115m@[0m[38;2;78;59;37mh[0m[38;2;76;61;43mh[0m[38;2;170;154;118m@[0m[38;2;177;160;121m@[0m[38;2;134;120;93mB[0m[38;2;52;40;23m2[0m[38;2;96;85;74mS[0m[38;2;42;32;18mX[0m[38;2;67;55;43mh[0m[38;2;58;47;35m5[0m[38;2;80;65;49mM[0m[38;2;103;90;71mS[0m[38;2;37;25;17ms[0m[38;2;126;114;86m9[0m[38;2;175;161;125m@[0m[38;2;174;159;121m@[0m[38;2;178;159;121m@[0m[38;2;163;138;104m&[0m[38;2;122;92;55mS[0m[38;2;124;92;52mS[0m[38;2;123;91;50mS[0m[38;2;124;90;50mS[0m[38;2;124;89;48mS[0m[38;2;145;108;66m9[0m[38;2;159;122;78mB[0m[38;2;160;123;78mB[0m[38;2;160;123;79mB[0m[38;2;161;123;79mB[0m[38;2;139;108;69m9[0m[38;2;91;67;35mM[0m[38;2;105;74;46mG[0m[38;2;129;93;60m#[0m[38;2;126;90;55m#[0m[38;2;131;92;57m#[0m[38;2;150;106;70m9[0m[38;2;157;112;77mB[0m[38;2;156;111;76mB[0m[38;2;159;115;79mB[0m[38;2;169;126;88m&[0m[38;2;176;133;95m&[0m[38;2;178;136;96m&[0m[38;2;177;136;95m&[0m[38;2;177;135;95m&[0m[38;2;177;135;95m&[0m[38;2;177;135;94m&[0m[38;2;177;135;94m&[0m[38;2;179;135;97m&[0m[38;2;178;135;95m&[0m[38;2;162;122;85mB[0m[38;2;130;89;64m#[0m[38;2;99;60;43mH[0m[38;2;89;53;36mh[0m[38;2;99;62;39mM[0m[38;2;115;77;49mG[0m[38;2;129;88;58m#[0m[38;2;119;82;51mS[0m[38;2;111;74;44mG[0m[38;2;115;78;50mG[0m[38;2;114;77;50mG[0m[38;2;109;72;47mG[0m[38;2;104;67;45mH[0m");
	$display("[38;2;90;62;42mM[0m[38;2;79;53;38mh[0m[38;2;73;48;37m3[0m[38;2;82;55;41mh[0m[38;2;101;72;53mG[0m[38;2;120;90;65m#[0m[38;2;145;110;79mB[0m[38;2;159;120;86mB[0m[38;2;164;121;87m&[0m[38;2;162;121;86mB[0m[38;2;163;123;88m&[0m[38;2;162;123;88m&[0m[38;2;163;123;88m&[0m[38;2;165;125;90m&[0m[38;2;165;126;91m&[0m[38;2;162;123;87m&[0m[38;2;154;115;79mB[0m[38;2;146;107;72m9[0m[38;2;149;110;72m9[0m[38;2;149;109;74mB[0m[38;2;136;97;68m9[0m[38;2;124;86;58mS[0m[38;2;136;98;68m9[0m[38;2;163;130;88m&[0m[38;2;140;108;68m9[0m[38;2;126;94;59m#[0m[38;2;124;91;58m#[0m[38;2;111;76;43mG[0m[38;2;142;106;66m9[0m[38;2;147;111;66m9[0m[38;2;149;111;68m9[0m[38;2;149;111;66m9[0m[38;2;148;112;65m9[0m[38;2;148;112;66m9[0m[38;2;148;112;66m9[0m[38;2;148;111;65m9[0m[38;2;147;111;65m9[0m[38;2;147;111;65m9[0m[38;2;146;111;65m9[0m[38;2;146;112;65m9[0m[38;2;145;111;64m9[0m[38;2;145;111;62m9[0m[38;2;158;130;87m&[0m[38;2;166;153;116m@[0m[38;2;71;59;46mh[0m[38;2;82;54;40mh[0m[38;2;194;153;114m@[0m[38;2;200;159;118m@[0m[38;2;192;156;113m@[0m[38;2;170;136;98m&[0m[38;2;152;118;90mB[0m[38;2;142;108;81m9[0m[38;2;150;116;85mB[0m[38;2;182;148;110m@[0m[38;2;194;162;114m@[0m[38;2;193;161;114m@[0m[38;2;194;161;116m@[0m[38;2;193;161;114m@[0m[38;2;193;161;115m@[0m[38;2;193;160;116m@[0m[38;2;193;160;117m@[0m[38;2;194;160;114m@[0m[38;2;194;161;112m@[0m[38;2;195;163;115m@[0m[38;2;187;157;115m@[0m[38;2;153;125;91mB[0m[38;2;126;98;70m#[0m[38;2;124;95;69m#[0m[38;2;128;99;70m#[0m[38;2;139;107;78m9[0m[38;2;153;123;91mB[0m[38;2;175;144;104m&[0m[38;2;193;157;113m@[0m[38;2;199;164;123m@[0m[38;2;133;108;78m9[0m[38;2;69;53;32m3[0m[38;2;165;150;115m@[0m[38;2;176;158;122m@[0m[38;2;118;103;81m9[0m[38;2;35;22;9mr[0m[38;2;58;46;36m5[0m[38;2;54;45;33m5[0m[38;2;32;24;15mr[0m[38;2;34;26;17ms[0m[38;2;41;29;20mX[0m[38;2;52;45;34m5[0m[38;2;31;25;20ms[0m[38;2;98;85;62mS[0m[38;2;176;157;124m@[0m[38;2;173;156;120m@[0m[38;2;174;157;122m@[0m[38;2;169;151;118m@[0m[38;2;123;98;62m#[0m[38;2;120;89;51mS[0m[38;2;122;90;50mS[0m[38;2;121;88;47mS[0m[38;2;122;86;45mS[0m[38;2;144;107;66m9[0m[38;2;159;122;78mB[0m[38;2;160;123;78mB[0m[38;2;161;123;79mB[0m[38;2;161;124;80mB[0m[38;2;140;110;70m9[0m[38;2;90;67;37mM[0m[38;2;97;67;43mH[0m[38;2;112;77;49mG[0m[38;2;129;90;60m#[0m[38;2;149;106;72m9[0m[38;2;155;110;72mB[0m[38;2;159;115;78mB[0m[38;2;167;126;89m&[0m[38;2;176;135;95m&[0m[38;2;177;136;96m&[0m[38;2;175;135;94m&[0m[38;2;174;135;93m&[0m[38;2;175;135;94m&[0m[38;2;176;134;95m&[0m[38;2;177;134;93m&[0m[38;2;176;134;93m&[0m[38;2;178;136;96m&[0m[38;2;168;127;92m&[0m[38;2;135;95;68m#[0m[38;2;97;59;40mM[0m[38;2;88;53;36mh[0m[38;2;95;62;43mM[0m[38;2;102;69;46mH[0m[38;2;109;73;48mG[0m[38;2;108;69;45mG[0m[38;2;110;72;50mG[0m[38;2;100;65;42mH[0m[38;2;94;61;39mM[0m[38;2;98;66;44mH[0m[38;2;99;66;42mH[0m[38;2;103;68;41mH[0m[38;2;112;75;44mG[0m");
	$display("[38;2;90;65;43mM[0m[38;2;96;67;45mH[0m[38;2;96;65;45mH[0m[38;2;86;58;43mM[0m[38;2;76;50;38mh[0m[38;2;69;45;34m3[0m[38;2;75;52;39mh[0m[38;2;105;76;59mG[0m[38;2;140;104;81m9[0m[38;2;158;118;87mB[0m[38;2;161;120;86mB[0m[38;2;162;121;86mB[0m[38;2;162;121;86mB[0m[38;2;162;123;87m&[0m[38;2;164;126;90m&[0m[38;2;165;127;91m&[0m[38;2;167;129;93m&[0m[38;2;164;126;90m&[0m[38;2;156;119;83mB[0m[38;2;149;110;74mB[0m[38;2;145;104;71m9[0m[38;2;137;97;68m9[0m[38;2;124;87;61m#[0m[38;2;121;87;58mS[0m[38;2;112;81;51mG[0m[38;2;117;89;58mS[0m[38;2;118;90;57mS[0m[38;2;108;76;42mG[0m[38;2;139;104;64m9[0m[38;2;145;109;63m9[0m[38;2;146;109;65m9[0m[38;2;147;110;64m9[0m[38;2;147;110;64m9[0m[38;2;146;109;65m9[0m[38;2;146;109;64m9[0m[38;2;146;109;64m9[0m[38;2;146;109;64m9[0m[38;2;146;109;64m9[0m[38;2;144;110;64m9[0m[38;2;144;110;64m9[0m[38;2;142;109;63m9[0m[38;2;142;110;62m9[0m[38;2;145;117;80mB[0m[38;2;163;148;116m&[0m[38;2;71;59;43mh[0m[38;2;82;58;41mh[0m[38;2;183;150;113m@[0m[38;2;161;131;96m&[0m[38;2;130;104;76m9[0m[38;2;119;96;70m#[0m[38;2;127;104;78m9[0m[38;2;122;102;73m#[0m[38;2;122;99;73m#[0m[38;2;139;112;82mB[0m[38;2;177;148;108m@[0m[38;2;191;159;114m@[0m[38;2;193;159;114m@[0m[38;2;193;160;115m@[0m[38;2;193;160;115m@[0m[38;2;193;160;115m@[0m[38;2;192;160;116m@[0m[38;2;193;159;115m@[0m[38;2;192;159;115m@[0m[38;2;169;139;99m&[0m[38;2;139;113;78m9[0m[38;2;134;110;78m9[0m[38;2;135;112;81m9[0m[38;2;141;118;87mB[0m[38;2;147;121;89mB[0m[38;2;141;115;83mB[0m[38;2;126;103;73m9[0m[38;2;115;96;68m#[0m[38;2;118;98;71m#[0m[38;2;138;114;86mB[0m[38;2;118;94;71m#[0m[38;2;68;53;36m3[0m[38;2;163;151;115m@[0m[38;2;173;158;119m@[0m[38;2;107;90;66mS[0m[38;2;59;46;34m5[0m[38;2;31;24;16mr[0m[38;2;31;25;12mr[0m[38;2;44;32;20mX[0m[38;2;53;42;27m2[0m[38;2;54;40;25m2[0m[38;2;37;27;17ms[0m[38;2;33;25;14mr[0m[38;2;74;61;43mh[0m[38;2;169;151;121m@[0m[38;2;170;154;116m@[0m[38;2;159;143;108m&[0m[38;2;171;156;121m@[0m[38;2;132;112;74m9[0m[38;2;117;87;49mS[0m[38;2;120;88;47mS[0m[38;2;119;88;44mS[0m[38;2;121;85;44mS[0m[38;2;143;105;64m9[0m[38;2;160;122;79mB[0m[38;2;161;123;79mB[0m[38;2;162;123;80mB[0m[38;2;162;124;81mB[0m[38;2;140;110;71m9[0m[38;2;87;62;36mM[0m[38;2;98;65;44mH[0m[38;2;125;89;61m#[0m[38;2;143;103;70m9[0m[38;2;157;113;78mB[0m[38;2;171;126;89m&[0m[38;2;176;134;96m&[0m[38;2;175;136;98m&[0m[38;2;174;136;96m&[0m[38;2;174;135;94m&[0m[38;2;174;135;94m&[0m[38;2;174;135;93m&[0m[38;2;175;134;94m&[0m[38;2;176;134;93m&[0m[38;2;176;134;92m&[0m[38;2;176;134;96m&[0m[38;2;151;111;80mB[0m[38;2;122;83;61mS[0m[38;2;102;64;45mH[0m[38;2;94;60;41mM[0m[38;2;99;68;47mH[0m[38;2;91;63;39mM[0m[38;2;82;54;31mh[0m[38;2;85;54;35mh[0m[38;2;91;58;40mM[0m[38;2;100;66;46mH[0m[38;2;99;65;42mH[0m[38;2;99;64;38mH[0m[38;2;117;81;49mS[0m[38;2;133;97;57m#[0m[38;2;149;112;67m9[0m[38;2;161;123;75mB[0m");
	$display("[38;2;65;45;27m5[0m[38;2;69;45;29m5[0m[38;2;79;51;34mh[0m[38;2;87;59;40mM[0m[38;2;92;65;44mH[0m[38;2;91;64;46mH[0m[38;2;82;58;42mM[0m[38;2;72;48;34m3[0m[38;2;74;49;34m3[0m[38;2;105;75;57mG[0m[38;2;143;108;84mB[0m[38;2;159;118;86mB[0m[38;2;159;118;82mB[0m[38;2;159;121;84mB[0m[38;2;160;123;87mB[0m[38;2;162;124;88m&[0m[38;2;163;126;90m&[0m[38;2;166;128;92m&[0m[38;2;166;128;93m&[0m[38;2;164;125;90m&[0m[38;2;157;117;82mB[0m[38;2;148;109;77mB[0m[38;2;138;102;72m9[0m[38;2;127;92;64m#[0m[38;2;103;71;46mH[0m[38;2;101;73;49mG[0m[38;2;105;79;51mG[0m[38;2;105;75;42mG[0m[38;2;139;104;60m9[0m[38;2;144;109;61m9[0m[38;2;145;108;64m9[0m[38;2;145;108;64m9[0m[38;2;145;108;64m9[0m[38;2;145;108;64m9[0m[38;2;144;108;63m9[0m[38;2;144;107;63m9[0m[38;2;144;107;63m9[0m[38;2;144;107;63m9[0m[38;2;142;108;63m9[0m[38;2;142;108;63m9[0m[38;2;140;107;61m9[0m[38;2;138;108;62m9[0m[38;2;139;113;77m9[0m[38;2;162;147;112m&[0m[38;2;72;63;45mh[0m[38;2;77;59;46mM[0m[38;2;122;98;71m#[0m[38;2;120;96;65m#[0m[38;2;153;127;92m&[0m[38;2;176;147;108m@[0m[38;2;186;153;111m@[0m[38;2;189;153;113m@[0m[38;2;184;150;111m@[0m[38;2;169;139;98m&[0m[38;2;174;146;103m&[0m[38;2;188;157;112m@[0m[38;2;192;158;113m@[0m[38;2;192;159;114m@[0m[38;2;191;158;113m@[0m[38;2;191;158;113m@[0m[38;2;191;159;115m@[0m[38;2;191;158;115m@[0m[38;2;189;156;116m@[0m[38;2;174;142;103m&[0m[38;2;178;145;107m@[0m[38;2;189;154;114m@[0m[38;2;192;159;115m@[0m[38;2;195;160;116m@[0m[38;2;196;156;115m@[0m[38;2;196;156;114m@[0m[38;2;192;154;112m@[0m[38;2;182;148;108m@[0m[38;2;164;134;98m&[0m[38;2;137;109;78m9[0m[38;2;88;68;47mH[0m[38;2;69;57;42mh[0m[38;2;165;151;119m@[0m[38;2;166;148;113m&[0m[38;2;101;80;58mG[0m[38;2;103;82;66mS[0m[38;2;64;43;24m5[0m[38;2;122;97;72m#[0m[38;2;138;104;84m9[0m[38;2;124;91;74m#[0m[38;2;112;87;63mS[0m[38;2;116;90;72m#[0m[38;2;49;30;19mX[0m[38;2;51;43;25m2[0m[38;2;155;140;111m&[0m[38;2;169;155;117m@[0m[38;2;155;140;103m&[0m[38;2;171;155;118m@[0m[38;2;146;127;90mB[0m[38;2;114;85;49mS[0m[38;2;118;86;47mS[0m[38;2;116;86;45mS[0m[38;2;119;84;44mS[0m[38;2;143;105;61m9[0m[38;2;158;121;76mB[0m[38;2;159;123;78mB[0m[38;2;158;123;80mB[0m[38;2;147;111;71m9[0m[38;2;120;88;53mS[0m[38;2;100;68;44mH[0m[38;2;124;83;60mS[0m[38;2;150;107;76mB[0m[38;2;167;123;88m&[0m[38;2;177;132;95m&[0m[38;2;176;134;95m&[0m[38;2;174;134;95m&[0m[38;2;174;134;98m&[0m[38;2;174;134;97m&[0m[38;2;173;134;95m&[0m[38;2;173;135;95m&[0m[38;2;174;135;94m&[0m[38;2;175;133;93m&[0m[38;2;174;134;95m&[0m[38;2;165;130;93m&[0m[38;2;126;92;65m#[0m[38;2;92;57;40mM[0m[38;2;95;61;46mH[0m[38;2;96;65;44mH[0m[38;2;92;63;38mM[0m[38;2;81;54;31mh[0m[38;2;77;50;29m3[0m[38;2;80;53;32mh[0m[38;2;92;61;38mM[0m[38;2;106;73;45mG[0m[38;2;133;98;63m#[0m[38;2;138;102;65m9[0m[38;2;141;104;62m9[0m[38;2;161;124;76mB[0m[38;2;167;128;76mB[0m[38;2;166;126;74mB[0m[38;2;164;126;74mB[0m");
	$display("[38;2;72;52;34m3[0m[38;2;67;48;32m3[0m[38;2;62;42;27m5[0m[38;2;60;38;24m2[0m[38;2;63;40;25m2[0m[38;2;71;47;31m3[0m[38;2;83;56;40mh[0m[38;2;91;64;50mH[0m[38;2;82;58;46mM[0m[38;2;71;48;35m3[0m[38;2;84;57;41mM[0m[38;2;118;85;64mS[0m[38;2;152;115;84mB[0m[38;2;159;119;83mB[0m[38;2;159;119;83mB[0m[38;2;159;120;84mB[0m[38;2;160;123;87mB[0m[38;2;163;124;88m&[0m[38;2;164;126;91m&[0m[38;2;165;127;91m&[0m[38;2;165;127;90m&[0m[38;2;163;125;89m&[0m[38;2;158;120;87mB[0m[38;2;150;112;82mB[0m[38;2;126;90;65m#[0m[38;2;107;74;53mG[0m[38;2;96;66;43mH[0m[38;2;99;69;40mH[0m[38;2;133;98;61m#[0m[38;2;143;107;63m9[0m[38;2;144;106;64m9[0m[38;2;142;106;64m9[0m[38;2;142;106;61m9[0m[38;2;142;106;61m9[0m[38;2;141;105;63m9[0m[38;2;140;105;62m9[0m[38;2;139;105;60m9[0m[38;2;140;105;60m9[0m[38;2;139;105;60m9[0m[38;2;139;105;60m9[0m[38;2;139;106;60m9[0m[38;2;137;105;61m9[0m[38;2;122;104;68m#[0m[38;2;159;146;112m&[0m[38;2;75;64;46mM[0m[38;2;60;43;28m5[0m[38;2;158;127;93m&[0m[38;2;188;148;108m@[0m[38;2;193;151;110m@[0m[38;2;191;149;110m@[0m[38;2;192;150;109m@[0m[38;2;192;154;113m@[0m[38;2;193;156;114m@[0m[38;2;194;158;116m@[0m[38;2;191;156;114m@[0m[38;2;192;158;116m@[0m[38;2;161;128;89m&[0m[38;2;156;122;86mB[0m[38;2;190;157;118m@[0m[38;2;190;157;114m@[0m[38;2;190;157;113m@[0m[38;2;190;157;114m@[0m[38;2;190;157;114m@[0m[38;2;192;158;115m@[0m[38;2;192;158;115m@[0m[38;2;190;156;114m@[0m[38;2;189;153;111m@[0m[38;2;189;149;108m@[0m[38;2;189;146;107m@[0m[38;2;191;145;108m@[0m[38;2;191;145;106m@[0m[38;2;193;149;108m@[0m[38;2;192;151;109m@[0m[38;2;194;153;114m@[0m[38;2;122;94;71m#[0m[38;2;78;64;45mM[0m[38;2;171;151;121m@[0m[38;2;147;130;104m&[0m[38;2;91;71;49mH[0m[38;2;112;85;63mS[0m[38;2;140;109;87mB[0m[38;2;100;73;59mG[0m[38;2;62;35;26m2[0m[38;2;45;24;19mX[0m[38;2;43;22;17ms[0m[38;2;112;78;66mS[0m[38;2;88;64;50mH[0m[38;2;33;28;13ms[0m[38;2;137;123;96mB[0m[38;2;173;156;119m@[0m[38;2;155;140;103m&[0m[38;2;169;152;117m@[0m[38;2;158;140;104m&[0m[38;2;112;88;51mS[0m[38;2;115;84;45mG[0m[38;2;116;83;43mG[0m[38;2;115;83;42mG[0m[38;2;133;101;61m#[0m[38;2;155;121;79mB[0m[38;2;147;113;69m9[0m[38;2;130;97;60m#[0m[38;2;120;86;59mS[0m[38;2;125;90;62m#[0m[38;2;137;101;67m9[0m[38;2;163;123;85mB[0m[38;2;174;132;95m&[0m[38;2;176;132;93m&[0m[38;2;175;133;93m&[0m[38;2;173;134;95m&[0m[38;2;172;133;95m&[0m[38;2;173;133;96m&[0m[38;2;173;132;94m&[0m[38;2;171;134;92m&[0m[38;2;171;134;93m&[0m[38;2;173;132;95m&[0m[38;2;173;132;97m&[0m[38;2;151;114;82mB[0m[38;2;110;76;50mG[0m[38;2;98;66;43mH[0m[38;2;106;74;51mG[0m[38;2;95;64;42mH[0m[38;2;86;56;34mh[0m[38;2;81;52;30m3[0m[38;2;82;55;32mh[0m[38;2;87;59;36mM[0m[38;2;99;67;42mH[0m[38;2;125;89;58m#[0m[38;2;145;106;68m9[0m[38;2;165;125;81mB[0m[38;2;160;123;77mB[0m[38;2;161;124;78mB[0m[38;2;170;132;84m&[0m[38;2;169;131;82m&[0m[38;2;167;128;78m&[0m[38;2;162;125;75mB[0m");
	$display("[38;2;117;90;52mS[0m[38;2;106;80;46mG[0m[38;2;94;69;41mH[0m[38;2;82;58;35mh[0m[38;2;72;50;30m3[0m[38;2;67;43;27m5[0m[38;2;62;39;24m2[0m[38;2;67;43;28m5[0m[38;2;79;53;38mh[0m[38;2;87;60;43mM[0m[38;2;80;56;40mh[0m[38;2;72;48;34m3[0m[38;2;96;65;48mH[0m[38;2;139;100;77m9[0m[38;2;157;117;85mB[0m[38;2;159;118;83mB[0m[38;2;159;119;83mB[0m[38;2;159;121;86mB[0m[38;2;160;121;87mB[0m[38;2;163;125;87m&[0m[38;2;165;126;87m&[0m[38;2;164;125;88m&[0m[38;2;164;125;90m&[0m[38;2;164;125;91m&[0m[38;2;159;119;89mB[0m[38;2;148;108;83mB[0m[38;2;122;87;62m#[0m[38;2;101;69;44mH[0m[38;2;107;75;46mG[0m[38;2;121;87;51mS[0m[38;2;135;99;62m#[0m[38;2;138;106;62m9[0m[38;2;136;105;59m9[0m[38;2;137;104;59m9[0m[38;2;139;103;59m9[0m[38;2;138;103;58m9[0m[38;2;136;104;58m#[0m[38;2;136;103;58m#[0m[38;2;136;103;58m#[0m[38;2;136;103;60m9[0m[38;2;136;103;60m9[0m[38;2;129;98;59m#[0m[38;2;97;82;51mG[0m[38;2;158;144;112m&[0m[38;2;81;69;53mH[0m[38;2;42;27;11ms[0m[38;2;161;123;93m&[0m[38;2;192;142;104m@[0m[38;2;192;140;101m@[0m[38;2;189;139;103m@[0m[38;2;192;142;104m@[0m[38;2;193;148;109m@[0m[38;2;193;154;112m@[0m[38;2;191;157;114m@[0m[38;2;189;156;113m@[0m[38;2;189;156;115m@[0m[38;2;175;142;103m&[0m[38;2;183;149;111m@[0m[38;2;189;156;116m@[0m[38;2;189;156;114m@[0m[38;2;189;156;113m@[0m[38;2;189;156;113m@[0m[38;2;189;156;113m@[0m[38;2;190;157;114m@[0m[38;2;190;156;113m@[0m[38;2;190;153;111m@[0m[38;2;189;147;107m@[0m[38;2;189;142;104m@[0m[38;2;190;140;102m@[0m[38;2;191;139;104m@[0m[38;2;190;139;102m@[0m[38;2;191;141;102m@[0m[38;2;190;140;103m@[0m[38;2;193;143;108m@[0m[38;2;114;83;62mS[0m[38;2;88;75;54mH[0m[38;2;172;154;123m@[0m[38;2;118;101;80m9[0m[38;2;103;78;49mG[0m[38;2;173;142;110m&[0m[38;2;95;67;50mH[0m[38;2;40;21;18ms[0m[38;2;43;27;24mX[0m[38;2;42;22;17ms[0m[38;2;53;25;19mX[0m[38;2;132;100;80m9[0m[38;2;84;64;45mM[0m[38;2;30;20;13mr[0m[38;2;116;100;80m#[0m[38;2;173;155;121m@[0m[38;2;155;140;106m&[0m[38;2;163;146;115m&[0m[38;2;168;150;118m@[0m[38;2;118;98;60m#[0m[38;2;111;85;43mG[0m[38;2;111;83;47mG[0m[38;2;103;77;49mG[0m[38;2;81;60;37mh[0m[38;2;91;68;49mH[0m[38;2;111;83;57mS[0m[38;2;126;90;57m#[0m[38;2;147;107;74m9[0m[38;2;164;125;88m&[0m[38;2;173;134;95m&[0m[38;2;173;134;94m&[0m[38;2;172;133;94m&[0m[38;2;172;133;94m&[0m[38;2;172;133;94m&[0m[38;2;172;133;94m&[0m[38;2;172;132;93m&[0m[38;2;172;131;91m&[0m[38;2;172;132;91m&[0m[38;2;173;132;91m&[0m[38;2;173;134;96m&[0m[38;2;164;125;92m&[0m[38;2;130;94;65m#[0m[38;2;105;69;44mH[0m[38;2;112;76;52mG[0m[38;2;116;80;56mS[0m[38;2;102;68;42mH[0m[38;2;83;55;30mh[0m[38;2;85;56;33mh[0m[38;2;95;66;42mH[0m[38;2;103;74;47mG[0m[38;2;107;78;48mG[0m[38;2;111;80;46mG[0m[38;2;132;95;59m#[0m[38;2;145;103;64m9[0m[38;2;151;109;66m9[0m[38;2;149;109;66m9[0m[38;2;147;108;65m9[0m[38;2;150;111;68m9[0m[38;2;160;121;77mB[0m[38;2;167;130;83m&[0m[38;2;168;130;82m&[0m");
	$display("[38;2;136;103;58m#[0m[38;2;136;103;59m#[0m[38;2;134;102;60m#[0m[38;2;130;98;58m#[0m[38;2;123;91;54mS[0m[38;2;110;81;47mG[0m[38;2;96;69;39mH[0m[38;2;80;56;32mh[0m[38;2;69;47;29m5[0m[38;2;65;44;28m5[0m[38;2;73;52;33m3[0m[38;2;84;61;39mM[0m[38;2;84;58;37mh[0m[38;2;84;56;38mh[0m[38;2;109;79;58mS[0m[38;2;143;109;82mB[0m[38;2;156;117;86mB[0m[38;2;159;116;82mB[0m[38;2;159;117;83mB[0m[38;2;159;120;86mB[0m[38;2;162;122;88m&[0m[38;2;164;124;91m&[0m[38;2;165;125;93m&[0m[38;2;165;125;91m&[0m[38;2;165;123;90m&[0m[38;2;167;124;92m&[0m[38;2;161;122;89m&[0m[38;2;145;109;77m9[0m[38;2;126;90;59m#[0m[38;2;112;77;49mG[0m[38;2;93;67;48mH[0m[38;2;82;61;40mM[0m[38;2;84;64;37mM[0m[38;2;107;83;51mG[0m[38;2;128;98;59m#[0m[38;2;137;103;60m9[0m[38;2;138;102;58m#[0m[38;2;134;101;57m#[0m[38;2;133;101;56m#[0m[38;2;133;101;58m#[0m[38;2;134;101;60m#[0m[38;2;127;94;60m#[0m[38;2;84;67;46mM[0m[38;2;153;136;111m&[0m[38;2;90;80;62mG[0m[38;2;26;19;8mi[0m[38;2;121;88;67m#[0m[38;2;189;142;107m@[0m[38;2;192;141;103m@[0m[38;2;189;143;107m@[0m[38;2;191;147;108m@[0m[38;2;191;152;111m@[0m[38;2;190;156;113m@[0m[38;2;189;157;113m@[0m[38;2;189;156;113m@[0m[38;2;189;156;113m@[0m[38;2;190;157;114m@[0m[38;2;190;157;112m@[0m[38;2;189;157;112m@[0m[38;2;189;157;112m@[0m[38;2;189;157;112m@[0m[38;2;189;156;113m@[0m[38;2;189;156;114m@[0m[38;2;189;156;115m@[0m[38;2;190;156;114m@[0m[38;2;190;154;113m@[0m[38;2;190;152;111m@[0m[38;2;191;150;109m@[0m[38;2;191;147;108m@[0m[38;2;190;146;107m@[0m[38;2;190;146;106m@[0m[38;2;190;145;105m@[0m[38;2;191;146;106m@[0m[38;2;192;148;112m@[0m[38;2;99;74;52mG[0m[38;2;100;89;66mS[0m[38;2;169;152;121m@[0m[38;2;86;67;51mH[0m[38;2;114;83;69mS[0m[38;2;129;98;82m9[0m[38;2;64;40;30m5[0m[38;2;40;21;16ms[0m[38;2;52;29;23mA[0m[38;2;89;60;43mM[0m[38;2;142;110;83mB[0m[38;2;124;98;75m#[0m[38;2;43;28;17mX[0m[38;2;30;20;14mr[0m[38;2;86;73;55mH[0m[38;2;169;152;120m@[0m[38;2;156;139;105m&[0m[38;2;150;132;104m&[0m[38;2;173;155;122m@[0m[38;2;135;114;82m9[0m[38;2;91;68;42mH[0m[38;2;85;64;41mM[0m[38;2;88;71;48mH[0m[38;2;60;48;33m5[0m[38;2;27;16;9mi[0m[38;2;68;46;33m3[0m[38;2;157;119;88mB[0m[38;2;174;131;91m&[0m[38;2;173;132;93m&[0m[38;2;172;131;94m&[0m[38;2;171;131;95m&[0m[38;2;170;132;96m&[0m[38;2;171;132;95m&[0m[38;2;171;132;94m&[0m[38;2;171;132;93m&[0m[38;2;172;131;92m&[0m[38;2;172;132;92m&[0m[38;2;173;132;94m&[0m[38;2;171;130;95m&[0m[38;2;146;106;77m9[0m[38;2;111;75;49mG[0m[38;2;105;72;49mG[0m[38;2;112;79;56mS[0m[38;2;107;74;51mG[0m[38;2;101;69;43mH[0m[38;2;107;76;48mG[0m[38;2;101;71;43mH[0m[38;2;105;75;49mG[0m[38;2;107;77;50mG[0m[38;2;107;77;47mG[0m[38;2;106;76;45mG[0m[38;2;107;76;45mG[0m[38;2;125;91;56m#[0m[38;2;137;100;60m#[0m[38;2;152;112;68mB[0m[38;2;159;118;73mB[0m[38;2;157;119;73mB[0m[38;2;149;113;68m9[0m[38;2;143;106;61m9[0m[38;2;147;110;65m9[0m[38;2;159;121;75mB[0m");
	$display("[38;2;133;100;59m#[0m[38;2;134;101;58m#[0m[38;2;134;101;58m#[0m[38;2;133;100;60m#[0m[38;2;134;100;61m#[0m[38;2;135;102;60m#[0m[38;2;134;101;59m#[0m[38;2;129;97;59m#[0m[38;2;116;87;53mS[0m[38;2;99;72;41mH[0m[38;2;79;54;30m3[0m[38;2;68;45;29m5[0m[38;2;73;49;36m3[0m[38;2;81;56;41mh[0m[38;2;82;54;38mh[0m[38;2;88;60;43mM[0m[38;2;118;86;65mS[0m[38;2;150;112;84mB[0m[38;2;160;118;86mB[0m[38;2;159;116;83mB[0m[38;2;159;118;84mB[0m[38;2;161;120;87mB[0m[38;2;162;122;90m&[0m[38;2;163;123;91m&[0m[38;2;165;125;92m&[0m[38;2;165;125;93m&[0m[38;2;164;125;92m&[0m[38;2;166;127;93m&[0m[38;2;157;122;93m&[0m[38;2;84;65;49mM[0m[38;2;21;15;9m;[0m[38;2;31;22;12mr[0m[38;2;65;50;38m3[0m[38;2;80;66;51mM[0m[38;2;84;68;45mM[0m[38;2;92;70;40mH[0m[38;2;118;90;57mS[0m[38;2;131;100;60m#[0m[38;2;132;100;56m#[0m[38;2;132;99;55m#[0m[38;2;133;99;58m#[0m[38;2;128;97;60m#[0m[38;2;81;67;45mM[0m[38;2;145;130;106m&[0m[38;2;100;91;68mS[0m[38;2;22;19;11mi[0m[38;2;72;51;34m3[0m[38;2;180;145;106m@[0m[38;2;191;152;109m@[0m[38;2;190;154;114m@[0m[38;2;189;155;110m@[0m[38;2;189;154;112m@[0m[38;2;189;155;112m@[0m[38;2;188;156;113m@[0m[38;2;189;156;113m@[0m[38;2;189;156;112m@[0m[38;2;192;159;115m@[0m[38;2;190;158;114m@[0m[38;2;190;157;112m@[0m[38;2;191;157;111m@[0m[38;2;192;157;114m@[0m[38;2;192;159;112m@[0m[38;2;193;160;114m@[0m[38;2;189;157;115m@[0m[38;2;188;155;116m@[0m[38;2;187;155;114m@[0m[38;2;186;156;113m@[0m[38;2;187;156;112m@[0m[38;2;190;155;113m@[0m[38;2;189;155;110m@[0m[38;2;190;154;111m@[0m[38;2;191;154;112m@[0m[38;2;190;154;112m@[0m[38;2;186;152;114m@[0m[38;2;83;65;42mM[0m[38;2;118;109;82m9[0m[38;2;153;136;107m&[0m[38;2;63;45;31m5[0m[38;2;108;81;67mS[0m[38;2;93;66;51mH[0m[38;2;97;69;49mH[0m[38;2;120;90;66m#[0m[38;2;135;104;79m9[0m[38;2;130;102;76m9[0m[38;2;84;63;51mM[0m[38;2;36;24;18ms[0m[38;2;32;22;13mr[0m[38;2;32;21;14mr[0m[38;2;57;46;32m5[0m[38;2;157;143;109m&[0m[38;2;161;145;107m&[0m[38;2;123;107;82m9[0m[38;2;140;124;103mB[0m[38;2;89;75;56mH[0m[38;2;52;42;29m2[0m[38;2;39;32;20mX[0m[38;2;48;39;25mA[0m[38;2;64;48;33m5[0m[38;2;54;45;28m2[0m[38;2;32;19;7mi[0m[38;2;117;86;68m#[0m[38;2;172;131;98m&[0m[38;2;171;131;94m&[0m[38;2;171;131;95m&[0m[38;2;171;131;95m&[0m[38;2;171;131;95m&[0m[38;2;171;131;96m&[0m[38;2;171;131;94m&[0m[38;2;171;132;92m&[0m[38;2;172;132;94m&[0m[38;2;172;131;97m&[0m[38;2;153;115;87mB[0m[38;2;120;84;61mS[0m[38;2;103;69;50mG[0m[38;2;105;72;52mG[0m[38;2;101;71;48mH[0m[38;2;99;68;43mH[0m[38;2;115;81;53mS[0m[38;2;140;105;71m9[0m[38;2;145;109;72m9[0m[38;2;112;79;47mG[0m[38;2;107;76;47mG[0m[38;2;104;75;47mG[0m[38;2;104;76;45mG[0m[38;2;104;74;43mH[0m[38;2;103;73;43mH[0m[38;2;118;86;53mS[0m[38;2;130;95;56m#[0m[38;2;147;109;63m9[0m[38;2;157;116;69mB[0m[38;2;156;118;71mB[0m[38;2;155;119;72mB[0m[38;2;154;118;72mB[0m[38;2;144;106;62m9[0m[38;2;139;100;57m#[0m");
	$display("[38;2;132;98;59m#[0m[38;2;132;99;58m#[0m[38;2;132;99;58m#[0m[38;2;132;98;60m#[0m[38;2;132;98;60m#[0m[38;2;133;99;58m#[0m[38;2;132;100;58m#[0m[38;2;133;100;58m#[0m[38;2;134;100;59m#[0m[38;2;136;99;60m#[0m[38;2;128;95;57m#[0m[38;2;108;83;48mG[0m[38;2;86;64;38mM[0m[38;2;68;45;27m5[0m[38;2;64;40;24m2[0m[38;2;66;45;33m5[0m[38;2;72;49;37m3[0m[38;2;92;61;45mM[0m[38;2;130;92;69m#[0m[38;2;153;113;84mB[0m[38;2;158;118;84mB[0m[38;2;157;117;83mB[0m[38;2;160;118;89mB[0m[38;2;159;120;88mB[0m[38;2;162;125;91m&[0m[38;2;162;127;92m&[0m[38;2;162;128;93m&[0m[38;2;160;127;95m&[0m[38;2;96;73;55mG[0m[38;2;27;19;10mi[0m[38;2;45;36;23mA[0m[38;2;50;38;28m2[0m[38;2;44;35;28mA[0m[38;2;25;21;15mr[0m[38;2;29;28;22ms[0m[38;2;44;39;26mA[0m[38;2;59;46;27m5[0m[38;2;84;65;40mM[0m[38;2;113;88;54mS[0m[38;2;130;98;57m#[0m[38;2;132;98;56m#[0m[38;2;130;99;60m#[0m[38;2;87;69;46mH[0m[38;2;126;109;85m9[0m[38;2;112;100;79m#[0m[38;2;26;19;14mi[0m[38;2;34;21;12mr[0m[38;2;130;105;74m9[0m[38;2;190;157;115m@[0m[38;2;186;155;113m@[0m[38;2;187;155;111m@[0m[38;2;189;154;111m@[0m[38;2;188;154;112m@[0m[38;2;188;155;112m@[0m[38;2;188;155;111m@[0m[38;2;173;138;105m&[0m[38;2;121;89;68m#[0m[38;2;130;104;85m9[0m[38;2;133;106;89m9[0m[38;2;132;103;84m9[0m[38;2;127;99;82m9[0m[38;2;104;79;64mS[0m[38;2;107;80;60mS[0m[38;2;171;139;104m&[0m[38;2;189;155;113m@[0m[38;2;188;155;114m@[0m[38;2;186;156;113m@[0m[38;2;187;156;112m@[0m[38;2;188;155;112m@[0m[38;2;188;155;110m@[0m[38;2;189;154;112m@[0m[38;2;190;154;112m@[0m[38;2;189;155;112m@[0m[38;2;178;146;109m@[0m[38;2;73;55;34m3[0m[38;2;139;129;100mB[0m[38;2;130;109;89m9[0m[38;2;60;36;27m2[0m[38;2;129;90;70m#[0m[38;2;147;108;85mB[0m[38;2;126;100;77m9[0m[38;2;77;63;46mM[0m[38;2;43;35;25mA[0m[38;2;26;22;16mr[0m[38;2;25;20;17mr[0m[38;2;28;24;14mr[0m[38;2;30;24;14mr[0m[38;2;31;21;18mr[0m[38;2;37;26;16ms[0m[38;2;130;116;95mB[0m[38;2;146;132;108m&[0m[38;2;78;66;49mM[0m[38;2;54;42;30m2[0m[38;2;37;28;19ms[0m[38;2;24;19;14mi[0m[38;2;17;13;8m;[0m[38;2;18;13;6m;[0m[38;2;54;42;31m2[0m[38;2;82;65;44mM[0m[38;2;43;30;20mX[0m[38;2;50;32;25mA[0m[38;2;155;121;95mB[0m[38;2;170;130;94m&[0m[38;2;170;130;94m&[0m[38;2;170;130;93m&[0m[38;2;170;131;92m&[0m[38;2;171;131;92m&[0m[38;2;171;132;90m&[0m[38;2;170;133;92m&[0m[38;2;161;124;92m&[0m[38;2;128;91;66m#[0m[38;2;103;68;47mH[0m[38;2;96;66;48mH[0m[38;2;90;64;44mM[0m[38;2;92;65;39mM[0m[38;2;112;83;48mG[0m[38;2;138;105;66m9[0m[38;2;154;117;76mB[0m[38;2;154;117;74mB[0m[38;2;143;110;67m9[0m[38;2;109;79;44mG[0m[38;2;103;76;44mG[0m[38;2;102;75;46mG[0m[38;2;103;73;45mH[0m[38;2;102;72;42mH[0m[38;2;103;70;39mH[0m[38;2;116;79;47mG[0m[38;2;125;84;50mS[0m[38;2;138;99;58m#[0m[38;2;149;107;64m9[0m[38;2;149;108;65m9[0m[38;2;148;109;65m9[0m[38;2;146;107;65m9[0m[38;2;145;105;63m9[0m[38;2;140;101;61m9[0m");
	$display("[38;2;131;97;59m#[0m[38;2;131;97;59m#[0m[38;2;131;97;59m#[0m[38;2;131;97;59m#[0m[38;2;132;98;60m#[0m[38;2;132;97;59m#[0m[38;2;132;97;59m#[0m[38;2;132;98;60m#[0m[38;2;132;98;60m#[0m[38;2;134;97;61m#[0m[38;2;132;97;58m#[0m[38;2;131;99;56m#[0m[38;2;128;98;59m#[0m[38;2;117;86;54mS[0m[38;2;93;66;39mM[0m[38;2;65;45;25m5[0m[38;2;53;36;21mA[0m[38;2;57;35;23m2[0m[38;2;70;43;29m5[0m[38;2;96;67;47mH[0m[38;2;133;99;73m9[0m[38;2;156;118;86mB[0m[38;2;160;118;85mB[0m[38;2;157;118;83mB[0m[38;2;157;121;86mB[0m[38;2;161;122;86mB[0m[38;2;160;125;91m&[0m[38;2;122;98;73m#[0m[38;2;48;38;22mA[0m[38;2;71;60;42mh[0m[38;2;88;73;45mH[0m[38;2;52;42;26m2[0m[38;2;19;15;10m;[0m[38;2;12;10;7m:[0m[38;2;10;10;8m:[0m[38;2;16;15;10m;[0m[38;2;30;26;18ms[0m[38;2;46;35;26mA[0m[38;2;59;45;31m5[0m[38;2;77;58;36mh[0m[38;2;105;79;49mG[0m[38;2;126;97;61m#[0m[38;2;105;83;55mG[0m[38;2;95;82;60mG[0m[38;2;117;106;85m9[0m[38;2;30;21;13mr[0m[38;2;26;20;14mr[0m[38;2;49;32;21mA[0m[38;2;150;121;91mB[0m[38;2;190;158;112m@[0m[38;2;188;156;109m@[0m[38;2;188;155;109m@[0m[38;2;188;155;110m@[0m[38;2;188;155;111m@[0m[38;2;188;155;113m@[0m[38;2;163;130;99m&[0m[38;2;45;20;13ms[0m[38;2;31;9;7mi[0m[38;2;54;25;20mX[0m[38;2;64;28;29m2[0m[38;2;64;28;27m2[0m[38;2;46;18;17ms[0m[38;2;58;31;22mA[0m[38;2;164;131;100m&[0m[38;2;191;154;112m@[0m[38;2;188;155;113m@[0m[38;2;188;155;113m@[0m[38;2;188;155;111m@[0m[38;2;188;155;111m@[0m[38;2;188;156;109m@[0m[38;2;189;154;114m@[0m[38;2;189;156;110m@[0m[38;2;190;160;112m@[0m[38;2;156;129;99m&[0m[38;2;74;59;38mh[0m[38;2;156;139;114m&[0m[38;2;90;76;59mG[0m[38;2;36;20;12mr[0m[38;2;51;27;21mX[0m[38;2;39;20;14ms[0m[38;2;24;21;12mi[0m[38;2;19;22;14mi[0m[38;2;23;23;18mr[0m[38;2;26;23;19mr[0m[38;2;27;23;18mr[0m[38;2;27;23;15mr[0m[38;2;36;33;23mX[0m[38;2;34;31;19ms[0m[38;2;31;21;11mr[0m[38;2;67;54;44mh[0m[38;2;62;50;41m3[0m[38;2;37;30;21mX[0m[38;2;22;17;10mi[0m[38;2;16;12;5m:[0m[38;2;16;13;6m;[0m[38;2;16;13;6m;[0m[38;2;14;13;5m:[0m[38;2;26;23;17mr[0m[38;2;37;27;19ms[0m[38;2;41;32;22mX[0m[38;2;23;10;9m;[0m[38;2;112;88;66mS[0m[38;2;168;131;93m&[0m[38;2;170;129;89m&[0m[38;2;168;130;93m&[0m[38;2;170;128;92m&[0m[38;2;171;130;95m&[0m[38;2;167;128;95m&[0m[38;2;143;107;78m9[0m[38;2;108;74;51mG[0m[38;2;96;65;44mH[0m[38;2;87;61;39mM[0m[38;2;83;60;37mh[0m[38;2;104;78;51mG[0m[38;2;133;102;67m9[0m[38;2;150;115;73mB[0m[38;2;153;115;72mB[0m[38;2;153;115;73mB[0m[38;2;152;115;73mB[0m[38;2;143;109;67m9[0m[38;2;106;78;44mG[0m[38;2;99;73;43mH[0m[38;2;100;72;45mH[0m[38;2;103;72;42mH[0m[38;2;111;78;44mG[0m[38;2;127;91;54m#[0m[38;2;136;97;61m#[0m[38;2;138;97;60m#[0m[38;2;137;98;58m#[0m[38;2;140;99;58m#[0m[38;2;140;99;57m#[0m[38;2;139;99;57m#[0m[38;2;138;98;56m#[0m[38;2;138;97;56m#[0m[38;2;139;98;59m#[0m");
	$display("[38;2;129;95;57m#[0m[38;2;129;95;57m#[0m[38;2;129;95;57m#[0m[38;2;129;96;57m#[0m[38;2;130;96;58m#[0m[38;2;130;96;58m#[0m[38;2;130;96;58m#[0m[38;2;130;96;58m#[0m[38;2;129;96;58m#[0m[38;2;130;96;58m#[0m[38;2;130;96;57m#[0m[38;2;130;96;55m#[0m[38;2;131;96;55m#[0m[38;2;131;97;56m#[0m[38;2;129;96;58m#[0m[38;2;118;90;55mS[0m[38;2;92;70;43mH[0m[38;2;62;43;25m5[0m[38;2;49;31;18mX[0m[38;2;54;34;23mA[0m[38;2;71;47;36m3[0m[38;2;104;71;55mG[0m[38;2;140;100;77m9[0m[38;2;157;117;84mB[0m[38;2;159;119;83mB[0m[38;2;161;117;82mB[0m[38;2;150;115;91mB[0m[38;2;54;39;28m2[0m[38;2;26;22;13mr[0m[38;2;48;37;26mA[0m[38;2;47;40;26mA[0m[38;2;31;26;19ms[0m[38;2;32;25;18ms[0m[38;2;29;24;17mr[0m[38;2;20;18;14mi[0m[38;2;13;12;9m:[0m[38;2;12;10;7m:[0m[38;2;17;12;9m;[0m[38;2;29;24;21ms[0m[38;2;37;32;28mX[0m[38;2;34;26;21ms[0m[38;2;53;41;27m2[0m[38;2;78;66;47mM[0m[38;2;72;62;42mh[0m[38;2;119;109;86m9[0m[38;2;28;24;15mr[0m[38;2;23;21;17mr[0m[38;2;29;23;15mr[0m[38;2;62;47;36m5[0m[38;2;122;95;71m#[0m[38;2;180;146;108m@[0m[38;2;191;157;116m@[0m[38;2;189;156;111m@[0m[38;2;187;155;109m@[0m[38;2;187;154;111m@[0m[38;2;189;154;116m@[0m[38;2;164;131;98m&[0m[38;2;143;101;76m9[0m[38;2;157;102;81mB[0m[38;2;162;103;85mB[0m[38;2;161;105;85mB[0m[38;2;166;117;90m&[0m[38;2;182;141;105m@[0m[38;2;189;153;113m@[0m[38;2;187;153;111m@[0m[38;2;187;155;112m@[0m[38;2;188;155;113m@[0m[38;2;189;155;112m@[0m[38;2;190;154;111m@[0m[38;2;192;156;113m@[0m[38;2;191;157;113m@[0m[38;2;182;150;109m@[0m[38;2;144;116;87mB[0m[38;2;73;52;34m3[0m[38;2;99;88;67mS[0m[38;2;134;119;96mB[0m[38;2;46;39;25mA[0m[38;2;23;21;16mr[0m[38;2;27;20;17mr[0m[38;2;28;21;17mr[0m[38;2;25;22;17mr[0m[38;2;26;23;17mr[0m[38;2;27;22;17mr[0m[38;2;26;22;15mr[0m[38;2;27;23;15mr[0m[38;2;25;21;12mi[0m[38;2;38;34;23mX[0m[38;2;53;49;37m5[0m[38;2;44;38;26mA[0m[38;2;35;28;21ms[0m[38;2;22;16;12mi[0m[38;2;17;12;8m;[0m[38;2;15;12;6m:[0m[38;2;16;13;6m;[0m[38;2;16;13;6m;[0m[38;2;16;12;6m:[0m[38;2;16;13;6m;[0m[38;2;14;11;7m:[0m[38;2;28;21;13mr[0m[38;2;36;32;19mX[0m[38;2;17;9;8m:[0m[38;2;66;47;31m5[0m[38;2;161;126;93m&[0m[38;2;170;129;86m&[0m[38;2;168;130;90m&[0m[38;2;170;130;96m&[0m[38;2;153;112;87mB[0m[38;2;118;83;61mS[0m[38;2;95;66;47mH[0m[38;2;87;60;42mM[0m[38;2;83;58;36mh[0m[38;2;96;73;43mH[0m[38;2;126;98;62m#[0m[38;2;146;112;72m9[0m[38;2;149;113;71mB[0m[38;2;148;112;69m9[0m[38;2;150;112;70mB[0m[38;2;150;112;72mB[0m[38;2;149;112;73mB[0m[38;2;141;107;69m9[0m[38;2;106;76;45mG[0m[38;2;99;70;42mH[0m[38;2;106;75;47mG[0m[38;2;124;90;57m#[0m[38;2;137;99;62m#[0m[38;2;141;102;63m9[0m[38;2;140;101;61m9[0m[38;2;140;101;61m9[0m[38;2;141;100;60m9[0m[38;2;140;101;61m9[0m[38;2;138;100;60m#[0m[38;2;138;100;60m#[0m[38;2;138;100;60m#[0m[38;2;138;100;60m#[0m[38;2;138;100;61m9[0m");
	$display("[38;2;126;95;55m#[0m[38;2;127;95;56m#[0m[38;2;127;95;56m#[0m[38;2;127;95;56m#[0m[38;2;127;95;56m#[0m[38;2;127;95;56m#[0m[38;2;127;96;56m#[0m[38;2;127;95;56m#[0m[38;2;127;95;56m#[0m[38;2;128;95;56m#[0m[38;2;128;95;56m#[0m[38;2;127;95;56m#[0m[38;2;127;96;56m#[0m[38;2;127;95;56m#[0m[38;2;128;95;55m#[0m[38;2;131;97;55m#[0m[38;2;125;93;55m#[0m[38;2;108;83;52mG[0m[38;2;85;64;40mM[0m[38;2;58;40;23m2[0m[38;2;46;29;19mX[0m[38;2;58;37;28m2[0m[38;2;77;51;38mh[0m[38;2;106;76;55mG[0m[38;2;143;105;76m9[0m[38;2;160;117;87mB[0m[38;2;114;87;70m#[0m[38;2;17;9;7m:[0m[38;2;23;19;15mi[0m[38;2;35;26;19ms[0m[38;2;13;12;7m:[0m[38;2;9;10;9m:[0m[38;2;17;12;7m;[0m[38;2;23;19;12mi[0m[38;2;28;25;17mr[0m[38;2;30;27;20ms[0m[38;2;27;23;18mr[0m[38;2;21;15;10m;[0m[38;2;14;10;5m:[0m[38;2;15;12;8m;[0m[38;2;25;21;16mr[0m[38;2;20;17;14mi[0m[38;2;25;23;20mr[0m[38;2;49;41;30m2[0m[38;2;118;105;87m9[0m[38;2;31;25;18ms[0m[38;2;23;19;16mi[0m[38;2;37;32;23mX[0m[38;2;54;52;40m5[0m[38;2;21;13;6m;[0m[38;2;68;47;36m3[0m[38;2;130;103;78m9[0m[38;2;175;142;105m&[0m[38;2;193;155;112m@[0m[38;2;192;156;114m@[0m[38;2;189;155;114m@[0m[38;2;189;157;110m@[0m[38;2;191;156;111m@[0m[38;2;189;153;113m@[0m[38;2;187;154;112m@[0m[38;2;188;155;112m@[0m[38;2;191;156;114m@[0m[38;2;189;155;113m@[0m[38;2;188;155;110m@[0m[38;2;187;155;110m@[0m[38;2;188;156;110m@[0m[38;2;192;158;109m@[0m[38;2;192;157;113m@[0m[38;2;185;149;113m@[0m[38;2;165;130;98m&[0m[38;2;123;94;70m#[0m[38;2;72;50;40m3[0m[38;2;32;18;12mr[0m[38;2;42;31;18mX[0m[38;2;130;117;99mB[0m[38;2;72;65;49mM[0m[38;2;27;25;16mr[0m[38;2;22;18;14mi[0m[38;2;30;25;21ms[0m[38;2;29;26;21ms[0m[38;2;25;23;16mr[0m[38;2;26;23;15mr[0m[38;2;25;21;13mi[0m[38;2;44;36;29mA[0m[38;2;37;28;22mX[0m[38;2;34;26;18ms[0m[38;2;43;35;27mA[0m[38;2;40;34;25mX[0m[38;2;24;20;11mi[0m[38;2;15;12;5m:[0m[38;2;14;12;7m:[0m[38;2;16;13;8m;[0m[38;2;16;13;7m;[0m[38;2;16;13;6m;[0m[38;2;16;13;6m;[0m[38;2;17;12;6m;[0m[38;2;16;12;6m:[0m[38;2;16;13;5m:[0m[38;2;46;39;26mA[0m[38;2;47;38;24mA[0m[38;2;25;16;12mi[0m[38;2;32;20;11mr[0m[38;2;141;111;84mB[0m[38;2;170;130;91m&[0m[38;2;156;119;85mB[0m[38;2;120;87;62mS[0m[38;2;94;63;44mH[0m[38;2;88;61;44mM[0m[38;2;81;56;38mh[0m[38;2;92;66;43mH[0m[38;2;120;91;62m#[0m[38;2;141;108;72m9[0m[38;2;147;112;73mB[0m[38;2;146;110;70m9[0m[38;2;144;111;71m9[0m[38;2;144;112;71m9[0m[38;2;144;111;70m9[0m[38;2;144;111;70m9[0m[38;2;144;111;70m9[0m[38;2;139;107;65m9[0m[38;2;113;79;40mG[0m[38;2;122;85;49mS[0m[38;2;136;97;63m#[0m[38;2;140;101;63m9[0m[38;2;141;100;61m9[0m[38;2;141;99;59m9[0m[38;2;140;100;59m9[0m[38;2;140;100;59m9[0m[38;2;141;100;60m9[0m[38;2;141;100;60m9[0m[38;2;141;100;61m9[0m[38;2;141;100;62m9[0m[38;2;140;99;61m9[0m[38;2;139;98;60m#[0m[38;2;138;100;59m#[0m");
	$display("[38;2;125;93;54m#[0m[38;2;125;93;54m#[0m[38;2;125;93;54m#[0m[38;2;126;94;55m#[0m[38;2;126;94;55m#[0m[38;2;125;93;54m#[0m[38;2;125;93;55m#[0m[38;2;125;93;54m#[0m[38;2;125;93;54m#[0m[38;2;126;94;55m#[0m[38;2;126;94;55m#[0m[38;2;126;94;55m#[0m[38;2;126;94;55m#[0m[38;2;126;94;55m#[0m[38;2;126;93;55m#[0m[38;2;128;93;54m#[0m[38;2;126;92;55m#[0m[38;2;114;83;49mS[0m[38;2;96;68;38mH[0m[38;2;86;61;35mM[0m[38;2;70;50;28m3[0m[38;2;53;35;19mA[0m[38;2;47;30;17mX[0m[38;2;57;40;27m2[0m[38;2;79;54;35mh[0m[38;2;105;78;58mG[0m[38;2;62;46;37m5[0m[38;2;11;6;5m,[0m[38;2;33;27;19ms[0m[38;2;47;41;30m2[0m[38;2;21;20;15mi[0m[38;2;10;9;7m:[0m[38;2;12;9;8m:[0m[38;2;14;11;7m:[0m[38;2;13;11;5m:[0m[38;2;18;15;9m;[0m[38;2;24;22;17mr[0m[38;2;31;28;23ms[0m[38;2;30;27;22ms[0m[38;2;23;20;15mi[0m[38;2;15;12;7m:[0m[38;2;16;12;7m;[0m[38;2;32;29;25mX[0m[38;2;34;26;17ms[0m[38;2;107;96;78m#[0m[38;2;32;27;18ms[0m[38;2;15;14;9m;[0m[38;2;39;30;25mX[0m[38;2;60;48;43m3[0m[38;2;22;15;13mi[0m[38;2;17;13;13m;[0m[38;2;22;16;13mi[0m[38;2;46;36;28mA[0m[38;2;87;69;53mH[0m[38;2;132;105;81m9[0m[38;2;170;137;103m&[0m[38;2;187;152;107m@[0m[38;2;193;156;112m@[0m[38;2;194;156;116m@[0m[38;2;192;157;113m@[0m[38;2;191;158;113m@[0m[38;2;191;158;114m@[0m[38;2;190;157;113m@[0m[38;2;187;154;111m@[0m[38;2;180;147;106m@[0m[38;2;165;133;98m&[0m[38;2;141;111;86mB[0m[38;2;111;83;68mS[0m[38;2;78;54;43mh[0m[38;2;51;30;23mA[0m[38;2;37;19;18ms[0m[38;2;30;18;18mr[0m[38;2;29;20;12mr[0m[38;2;89;81;63mG[0m[38;2;84;74;54mH[0m[38;2;35;30;19ms[0m[38;2;18;16;11m;[0m[38;2;10;4;3m,[0m[38;2;38;29;27mX[0m[38;2;38;30;27mX[0m[38;2;25;21;15mr[0m[38;2;24;21;15mr[0m[38;2;25;21;14mr[0m[38;2;55;46;37m5[0m[38;2;50;42;33m2[0m[38;2;37;32;25mX[0m[38;2;25;22;16mr[0m[38;2;14;12;8m:[0m[38;2;14;11;7m:[0m[38;2;14;12;7m:[0m[38;2;14;12;7m:[0m[38;2;15;12;7m:[0m[38;2;15;12;7m:[0m[38;2;15;12;7m:[0m[38;2;15;12;7m:[0m[38;2;15;12;7m:[0m[38;2;15;12;8m;[0m[38;2;13;11;7m:[0m[38;2;32;28;19ms[0m[38;2;48;35;26mA[0m[38;2;40;30;23mX[0m[38;2;18;10;4m:[0m[38;2;104;81;65mS[0m[38;2;125;91;69m#[0m[38;2;81;50;32m3[0m[38;2;75;50;34m3[0m[38;2;77;54;35mh[0m[38;2;84;59;36mh[0m[38;2;113;83;55mS[0m[38;2;139;105;70m9[0m[38;2;146;109;71m9[0m[38;2;145;108;68m9[0m[38;2;145;108;69m9[0m[38;2;145;108;69m9[0m[38;2;145;107;68m9[0m[38;2;144;107;68m9[0m[38;2;144;108;68m9[0m[38;2;144;108;68m9[0m[38;2;144;108;68m9[0m[38;2;145;108;69m9[0m[38;2;143;107;67m9[0m[38;2;149;109;69m9[0m[38;2;151;109;66m9[0m[38;2;150;109;64m9[0m[38;2;149;110;64m9[0m[38;2;148;110;65m9[0m[38;2;149;110;65m9[0m[38;2;149;111;66m9[0m[38;2;149;111;66m9[0m[38;2;148;109;64m9[0m[38;2;146;108;63m9[0m[38;2;147;108;64m9[0m[38;2;146;107;64m9[0m[38;2;146;106;64m9[0m[38;2;147;106;63m9[0m");
	$display("[38;2;124;92;54m#[0m[38;2;124;92;54m#[0m[38;2;124;92;54m#[0m[38;2;124;92;54m#[0m[38;2;124;92;54m#[0m[38;2;124;92;54m#[0m[38;2;125;93;55m#[0m[38;2;124;92;54m#[0m[38;2;124;92;54m#[0m[38;2;124;92;54m#[0m[38;2;124;92;54m#[0m[38;2;124;92;54m#[0m[38;2;124;92;54m#[0m[38;2;124;92;54m#[0m[38;2;124;92;54m#[0m[38;2;123;92;54mS[0m[38;2;123;92;54mS[0m[38;2;121;92;53mS[0m[38;2;119;87;50mS[0m[38;2;118;86;50mS[0m[38;2;113;85;49mS[0m[38;2;93;69;39mH[0m[38;2;72;51;28m3[0m[38;2;61;40;21m2[0m[38;2;55;34;18mA[0m[38;2;57;41;30m2[0m[38;2;23;16;11mi[0m[38;2;23;18;15mi[0m[38;2;46;35;28mA[0m[38;2;34;27;21ms[0m[38;2;13;13;12m;[0m[38;2;11;9;9m:[0m[38;2;12;9;9m:[0m[38;2;12;10;10m:[0m[38;2;12;11;7m:[0m[38;2;12;11;7m:[0m[38;2;12;11;9m:[0m[38;2;14;13;10m;[0m[38;2;19;18;15mi[0m[38;2;28;27;23ms[0m[38;2;28;27;22ms[0m[38;2;14;12;5m:[0m[38;2;27;25;20mr[0m[38;2;26;20;13mi[0m[38;2;80;68;54mH[0m[38;2;47;34;26mA[0m[38;2;25;12;10mi[0m[38;2;19;11;9m;[0m[38;2;37;27;26mX[0m[38;2;36;24;24ms[0m[38;2;9;6;4m,[0m[38;2;5;3;1m.[0m[38;2;1;2;2m.[0m[38;2;0;0;0m [0m[38;2;2;1;1m.[0m[38;2;34;26;21ms[0m[38;2;73;58;43mh[0m[38;2;109;87;65mS[0m[38;2;139;109;85mB[0m[38;2;150;117;87mB[0m[38;2;144;112;82mB[0m[38;2;131;101;75m9[0m[38;2;111;83;64mS[0m[38;2;89;64;51mH[0m[38;2;67;45;35m3[0m[38;2;51;30;24mA[0m[38;2;39;21;19ms[0m[38;2;35;19;18mr[0m[38;2;36;21;18ms[0m[38;2;38;23;18ms[0m[38;2;38;24;19ms[0m[38;2;32;21;17mr[0m[38;2;55;47;41m5[0m[38;2;61;55;47m3[0m[38;2;34;29;21ms[0m[38;2;19;18;14mi[0m[38;2;4;3;4m.[0m[38;2;8;5;5m,[0m[38;2;41;36;33mA[0m[38;2;34;28;25mX[0m[38;2;24;21;15mr[0m[38;2;33;32;24mX[0m[38;2;40;36;29mA[0m[38;2;32;28;21ms[0m[38;2;22;17;12mi[0m[38;2;14;11;8m:[0m[38;2;12;11;8m:[0m[38;2;12;11;10m:[0m[38;2;12;11;8m:[0m[38;2;12;11;8m:[0m[38;2;12;11;8m:[0m[38;2;12;12;7m:[0m[38;2;13;11;8m:[0m[38;2;13;11;9m:[0m[38;2;13;11;9m:[0m[38;2;13;11;8m:[0m[38;2;12;11;8m:[0m[38;2;11;11;7m:[0m[38;2;14;13;7m:[0m[38;2;45;36;28mA[0m[38;2;56;45;35m5[0m[38;2;26;22;12mr[0m[38;2;36;27;19ms[0m[38;2;52;34;25mA[0m[38;2;42;23;16ms[0m[38;2;60;36;25m2[0m[38;2;94;64;41mM[0m[38;2;126;93;64m#[0m[38;2;142;107;71m9[0m[38;2;143;107;68m9[0m[38;2;142;107;67m9[0m[38;2;142;107;68m9[0m[38;2;141;106;68m9[0m[38;2;142;106;68m9[0m[38;2;141;106;68m9[0m[38;2;141;106;67m9[0m[38;2;143;107;69m9[0m[38;2;143;107;69m9[0m[38;2;143;107;69m9[0m[38;2;143;107;69m9[0m[38;2;144;108;68m9[0m[38;2;146;109;67m9[0m[38;2;147;109;66m9[0m[38;2;145;109;65m9[0m[38;2;145;110;65m9[0m[38;2;146;109;65m9[0m[38;2;145;108;64m9[0m[38;2;145;108;64m9[0m[38;2;145;108;64m9[0m[38;2;144;107;65m9[0m[38;2;144;106;65m9[0m[38;2;143;105;65m9[0m[38;2;142;104;65m9[0m[38;2;142;104;65m9[0m[38;2;141;104;63m9[0m");
	$display("[38;2;123;91;53mS[0m[38;2;123;91;53mS[0m[38;2;123;91;53mS[0m[38;2;123;91;53mS[0m[38;2;123;91;53mS[0m[38;2;123;91;53mS[0m[38;2;123;91;53mS[0m[38;2;124;91;53mS[0m[38;2;124;92;54m#[0m[38;2;122;92;54mS[0m[38;2;122;92;54mS[0m[38;2;122;92;54mS[0m[38;2;122;92;54mS[0m[38;2;121;91;53mS[0m[38;2;121;91;53mS[0m[38;2;121;91;53mS[0m[38;2;120;91;53mS[0m[38;2;121;91;53mS[0m[38;2;122;91;54mS[0m[38;2;123;92;53mS[0m[38;2;117;88;50mS[0m[38;2;97;72;39mH[0m[38;2;87;63;37mM[0m[38;2;96;71;47mH[0m[38;2;80;55;32mh[0m[38;2;52;36;23mA[0m[38;2;17;12;5m:[0m[38;2;45;38;26mA[0m[38;2;61;49;35m5[0m[38;2;31;26;18ms[0m[38;2;12;11;8m:[0m[38;2;12;11;7m:[0m[38;2;10;11;8m:[0m[38;2;11;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;8m:[0m[38;2;11;12;7m:[0m[38;2;12;11;8m:[0m[38;2;12;11;9m:[0m[38;2;14;13;10m;[0m[38;2;20;19;14mi[0m[38;2;18;18;10m;[0m[38;2;22;22;17mr[0m[38;2;26;24;20mr[0m[38;2;39;30;24mX[0m[38;2;63;46;36m5[0m[38;2;105;67;59mG[0m[38;2;60;23;22mA[0m[38;2;18;10;9m;[0m[38;2;11;5;6m,[0m[38;2;4;4;3m.[0m[38;2;0;1;1m.[0m[38;2;0;0;0m [0m[38;2;0;0;0m [0m[38;2;0;0;1m.[0m[38;2;0;1;2m.[0m[38;2;12;11;9m:[0m[38;2;21;15;9m;[0m[38;2;28;16;12mi[0m[38;2;39;23;23ms[0m[38;2;38;22;20ms[0m[38;2;38;19;18ms[0m[38;2;37;18;17mr[0m[38;2;35;20;17mr[0m[38;2;34;22;19ms[0m[38;2;37;23;21ms[0m[38;2;38;24;21ms[0m[38;2;39;24;21ms[0m[38;2;39;24;21ms[0m[38;2;38;23;21ms[0m[38;2;34;22;19ms[0m[38;2;30;21;17mr[0m[38;2;31;26;21ms[0m[38;2;27;24;18mr[0m[38;2;17;16;12m;[0m[38;2;4;3;2m.[0m[38;2;1;0;0m.[0m[38;2;5;4;3m,[0m[38;2;16;14;13m;[0m[38;2;14;9;8m:[0m[38;2;29;27;21ms[0m[38;2;38;40;30mA[0m[38;2;23;18;11mi[0m[38;2;13;9;7m:[0m[38;2;13;9;8m:[0m[38;2;13;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;8m:[0m[38;2;12;11;7m:[0m[38;2;50;40;29m2[0m[38;2;76;61;44mh[0m[38;2;38;30;18mX[0m[38;2;20;13;12m;[0m[38;2;34;24;17ms[0m[38;2;20;8;6m:[0m[38;2;60;39;30m2[0m[38;2;117;82;59mS[0m[38;2;133;97;67m#[0m[38;2;139;105;67m9[0m[38;2;139;106;65m9[0m[38;2;138;105;65m9[0m[38;2;139;105;67m9[0m[38;2;140;106;68m9[0m[38;2;139;106;68m9[0m[38;2;138;104;66m9[0m[38;2;139;104;66m9[0m[38;2;139;104;66m9[0m[38;2;140;105;67m9[0m[38;2;139;105;67m9[0m[38;2;139;104;66m9[0m[38;2;141;104;66m9[0m[38;2;143;106;65m9[0m[38;2;143;106;63m9[0m[38;2;144;107;65m9[0m[38;2;144;107;65m9[0m[38;2;143;106;64m9[0m[38;2;143;106;64m9[0m[38;2;143;106;63m9[0m[38;2;142;105;62m9[0m[38;2;142;104;65m9[0m[38;2;142;104;65m9[0m[38;2;141;103;64m9[0m[38;2;139;101;62m9[0m[38;2;140;102;63m9[0m[38;2;140;102;63m9[0m");
	$display("[38;2;122;89;52mS[0m[38;2;122;90;52mS[0m[38;2;122;90;52mS[0m[38;2;122;89;52mS[0m[38;2;121;89;52mS[0m[38;2;120;89;52mS[0m[38;2;120;90;52mS[0m[38;2;121;90;52mS[0m[38;2;120;90;52mS[0m[38;2;120;90;52mS[0m[38;2;120;90;52mS[0m[38;2;120;90;52mS[0m[38;2;120;90;52mS[0m[38;2;120;90;52mS[0m[38;2;120;90;52mS[0m[38;2;120;90;52mS[0m[38;2;120;90;52mS[0m[38;2;120;90;52mS[0m[38;2;121;90;53mS[0m[38;2;122;90;52mS[0m[38;2;116;89;51mS[0m[38;2;99;74;41mH[0m[38;2;85;61;35mh[0m[38;2;96;71;45mH[0m[38;2;95;69;40mH[0m[38;2;76;59;38mh[0m[38;2;28;20;8mi[0m[38;2;60;51;36m3[0m[38;2;79;66;47mM[0m[38;2;44;35;25mA[0m[38;2;23;19;13mi[0m[38;2;17;17;11m;[0m[38;2;14;16;10m;[0m[38;2;16;16;12m;[0m[38;2;18;16;11m;[0m[38;2;19;17;11mi[0m[38;2;17;17;10m;[0m[38;2;14;14;8m;[0m[38;2;13;12;8m:[0m[38;2;12;11;8m:[0m[38;2;13;13;8m:[0m[38;2;20;17;11mi[0m[38;2;24;16;11mi[0m[38;2;39;31;24mX[0m[38;2;49;41;31m2[0m[38;2;31;21;9mr[0m[38;2;58;14;13ms[0m[38;2;58;3;9mr[0m[38;2;13;1;0m,[0m[38;2;4;4;3m.[0m[38;2;11;11;12m:[0m[38;2;8;8;8m:[0m[38;2;2;2;2m.[0m[38;2;1;1;1m.[0m[38;2;1;1;1m.[0m[38;2;0;1;0m.[0m[38;2;2;2;1m.[0m[38;2;16;12;9m;[0m[38;2;27;17;15mi[0m[38;2;36;23;23ms[0m[38;2;36;24;21ms[0m[38;2;38;24;21ms[0m[38;2;39;24;21ms[0m[38;2;39;24;20ms[0m[38;2;39;24;20ms[0m[38;2;39;24;21ms[0m[38;2;39;24;21ms[0m[38;2;39;24;21ms[0m[38;2;39;24;21ms[0m[38;2;37;22;19ms[0m[38;2;35;22;20ms[0m[38;2;30;20;19mr[0m[38;2;24;18;16mi[0m[38;2;21;17;14mi[0m[38;2;5;4;1m.[0m[38;2;1;0;0m.[0m[38;2;6;4;5m,[0m[38;2;12;11;10m:[0m[38;2;10;8;8m:[0m[38;2;8;8;6m,[0m[38;2;15;13;9m;[0m[38;2;23;16;13mi[0m[38;2;12;10;7m:[0m[38;2;14;10;9m:[0m[38;2;14;10;9m:[0m[38;2;13;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;8m:[0m[38;2;12;11;8m:[0m[38;2;11;11;7m:[0m[38;2;34;26;17ms[0m[38;2;49;37;24mA[0m[38;2;32;26;16ms[0m[38;2;14;8;11m:[0m[38;2;10;6;4m,[0m[38;2;5;0;0m.[0m[38;2;60;43;32m5[0m[38;2;113;79;54mS[0m[38;2;130;94;63m#[0m[38;2;136;102;65m9[0m[38;2;137;104;65m9[0m[38;2;136;102;65m9[0m[38;2;136;102;64m9[0m[38;2;135;101;63m9[0m[38;2;135;101;63m9[0m[38;2;135;101;64m9[0m[38;2;135;101;63m9[0m[38;2;135;101;63m9[0m[38;2;136;101;63m9[0m[38;2;136;102;64m9[0m[38;2;137;103;65m9[0m[38;2;139;102;65m9[0m[38;2;140;104;63m9[0m[38;2;140;104;61m9[0m[38;2;140;104;62m9[0m[38;2;141;104;64m9[0m[38;2;141;103;63m9[0m[38;2;140;103;62m9[0m[38;2;140;103;62m9[0m[38;2;139;102;61m9[0m[38;2;139;101;62m9[0m[38;2;139;101;62m9[0m[38;2;138;100;61m9[0m[38;2;136;98;59m#[0m[38;2;138;99;60m#[0m[38;2;139;101;62m9[0m");
	$display("[38;2;119;89;50mS[0m[38;2;119;89;49mS[0m[38;2;119;89;49mS[0m[38;2;119;89;50mS[0m[38;2;118;89;50mS[0m[38;2;118;89;50mS[0m[38;2;118;89;49mS[0m[38;2;118;89;50mS[0m[38;2;119;89;50mS[0m[38;2;120;89;50mS[0m[38;2;120;89;50mS[0m[38;2;120;89;50mS[0m[38;2;120;89;50mS[0m[38;2;120;89;50mS[0m[38;2;119;89;50mS[0m[38;2;118;89;49mS[0m[38;2;118;89;50mS[0m[38;2;118;89;49mS[0m[38;2;118;88;51mS[0m[38;2;119;88;50mS[0m[38;2;118;87;50mS[0m[38;2;103;77;45mG[0m[38;2;84;62;36mM[0m[38;2;92;68;41mH[0m[38;2;87;61;33mh[0m[38;2;71;53;32m3[0m[38;2;44;32;21mX[0m[38;2;57;47;35m5[0m[38;2;57;46;31m5[0m[38;2;47;36;26mA[0m[38;2;40;32;25mX[0m[38;2;29;25;18mr[0m[38;2;25;24;17mr[0m[38;2;28;25;19mr[0m[38;2;34;28;21ms[0m[38;2;37;30;22mX[0m[38;2;38;33;24mX[0m[38;2;36;31;24mX[0m[38;2;29;23;19mr[0m[38;2;19;15;12m;[0m[38;2;20;14;11m;[0m[38;2;35;9;7mi[0m[38;2;64;29;24m2[0m[38;2;55;28;21mA[0m[38;2;57;27;21mA[0m[38;2;40;13;8mr[0m[38;2;44;12;12mr[0m[38;2;59;7;15ms[0m[38;2;34;5;8mi[0m[38;2;12;9;6m:[0m[38;2;12;9;8m:[0m[38;2;10;10;9m:[0m[38;2;3;3;2m.[0m[38;2;1;1;1m.[0m[38;2;1;1;1m.[0m[38;2;1;1;1m.[0m[38;2;1;0;1m.[0m[38;2;5;0;1m.[0m[38;2;26;15;14mi[0m[38;2;39;22;20ms[0m[38;2;37;22;18ms[0m[38;2;37;23;19ms[0m[38;2;38;23;20ms[0m[38;2;39;22;20ms[0m[38;2;39;22;20ms[0m[38;2;38;23;20ms[0m[38;2;39;24;21ms[0m[38;2;39;24;21ms[0m[38;2;39;24;21ms[0m[38;2;39;24;21ms[0m[38;2;39;23;22ms[0m[38;2;36;22;21ms[0m[38;2;22;15;13mi[0m[38;2;8;7;5m,[0m[38;2;4;3;3m.[0m[38;2;11;10;10m:[0m[38;2;18;16;16mi[0m[38;2;15;12;12m;[0m[38;2;4;2;1m.[0m[38;2;1;3;1m.[0m[38;2;19;4;3m:[0m[38;2;38;4;7mi[0m[38;2;19;9;9m;[0m[38;2;11;12;8m:[0m[38;2;13;11;8m:[0m[38;2;12;11;8m:[0m[38;2;12;11;9m:[0m[38;2;14;10;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;12;11;9m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;12;10;8m:[0m[38;2;15;11;3m:[0m[38;2;31;28;20ms[0m[38;2;23;22;18mr[0m[38;2;10;7;8m:[0m[38;2;4;1;2m.[0m[38;2;8;1;1m.[0m[38;2;67;47;36m3[0m[38;2;108;76;49mG[0m[38;2;126;92;57m#[0m[38;2;134;98;63m#[0m[38;2;136;100;66m9[0m[38;2;133;99;62m#[0m[38;2;132;98;60m#[0m[38;2;132;98;60m#[0m[38;2;132;98;61m#[0m[38;2;132;98;61m#[0m[38;2;132;98;60m#[0m[38;2;133;99;62m#[0m[38;2;134;100;62m#[0m[38;2;134;100;62m#[0m[38;2;134;100;62m#[0m[38;2;135;100;63m#[0m[38;2;137;102;64m9[0m[38;2;137;102;64m9[0m[38;2;137;102;64m9[0m[38;2;137;102;64m9[0m[38;2;137;101;64m9[0m[38;2;137;100;63m9[0m[38;2;138;99;63m9[0m[38;2;137;99;62m#[0m[38;2;137;99;61m#[0m[38;2;137;98;61m#[0m[38;2;137;99;61m#[0m[38;2;137;98;59m#[0m[38;2;137;98;59m#[0m[38;2;137;98;59m#[0m");
	$display("[38;2;117;88;49mS[0m[38;2;117;87;49mS[0m[38;2;117;87;49mS[0m[38;2;117;88;49mS[0m[38;2;117;87;49mS[0m[38;2;118;88;49mS[0m[38;2;117;87;49mS[0m[38;2;117;87;49mS[0m[38;2;117;87;49mS[0m[38;2;118;87;49mS[0m[38;2;118;87;49mS[0m[38;2;118;87;49mS[0m[38;2;118;88;49mS[0m[38;2;118;87;49mS[0m[38;2;117;87;49mS[0m[38;2;117;87;49mS[0m[38;2;117;87;49mS[0m[38;2;117;87;49mS[0m[38;2;117;87;50mS[0m[38;2;118;87;49mS[0m[38;2;118;86;49mS[0m[38;2;105;79;46mG[0m[38;2;86;65;39mM[0m[38;2;90;67;42mM[0m[38;2;84;57;31mh[0m[38;2;75;56;36mh[0m[38;2;44;34;23mA[0m[38;2;45;36;25mA[0m[38;2;52;43;29m2[0m[38;2;51;41;30m2[0m[38;2;35;27;18ms[0m[38;2;27;24;17mr[0m[38;2;24;21;15mr[0m[38;2;25;20;15mr[0m[38;2;29;21;17mr[0m[38;2;31;23;20ms[0m[38;2;32;25;20ms[0m[38;2;33;25;21ms[0m[38;2;28;24;21ms[0m[38;2;23;18;14mi[0m[38;2;39;8;8mi[0m[38;2;71;21;17mA[0m[38;2;137;94;80m9[0m[38;2;65;30;20m2[0m[38;2;53;10;8mr[0m[38;2;62;8;12ms[0m[38;2;48;9;13mr[0m[38;2;30;9;11mi[0m[38;2;15;10;10m;[0m[38;2;10;10;10m:[0m[38;2;11;9;9m:[0m[38;2;11;11;9m:[0m[38;2;4;4;3m.[0m[38;2;1;1;1m.[0m[38;2;1;1;1m.[0m[38;2;1;1;1m.[0m[38;2;2;1;1m.[0m[38;2;4;0;1m.[0m[38;2;26;14;14mi[0m[38;2;38;20;19ms[0m[38;2;35;19;16mr[0m[38;2;35;20;17mr[0m[38;2;35;19;17mr[0m[38;2;36;20;19ms[0m[38;2;36;20;19ms[0m[38;2;37;22;20ms[0m[38;2;37;22;19ms[0m[38;2;37;22;19ms[0m[38;2;37;22;19ms[0m[38;2;38;22;21ms[0m[38;2;40;23;23mX[0m[38;2;29;15;15mi[0m[38;2;10;3;2m,[0m[38;2;10;9;6m:[0m[38;2;13;15;10m;[0m[38;2;13;13;9m;[0m[38;2;13;10;7m:[0m[38;2;14;8;6m:[0m[38;2;18;3;5m:[0m[38;2;31;7;7m;[0m[38;2;105;67;57mG[0m[38;2;91;41;32mh[0m[38;2;45;2;5mi[0m[38;2;19;9;6m:[0m[38;2;10;11;6m:[0m[38;2;12;10;9m:[0m[38;2;12;9;9m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;10;10;8m:[0m[38;2;16;11;11m;[0m[38;2;44;39;30mA[0m[38;2;35;30;21mX[0m[38;2;14;11;9m:[0m[38;2;11;6;6m:[0m[38;2;4;0;1m.[0m[38;2;11;4;2m,[0m[38;2;74;55;40mh[0m[38;2;106;75;46mG[0m[38;2;123;90;53mS[0m[38;2;132;97;60m#[0m[38;2;132;97;62m#[0m[38;2;130;97;59m#[0m[38;2;129;95;58m#[0m[38;2;129;95;58m#[0m[38;2;131;97;60m#[0m[38;2;130;96;59m#[0m[38;2;130;96;59m#[0m[38;2;131;97;60m#[0m[38;2;130;96;59m#[0m[38;2;131;97;59m#[0m[38;2;132;98;60m#[0m[38;2;133;99;61m#[0m[38;2;134;100;62m#[0m[38;2;134;100;62m#[0m[38;2;134;99;61m#[0m[38;2;134;99;61m#[0m[38;2;134;99;61m#[0m[38;2;135;98;61m#[0m[38;2;136;98;61m#[0m[38;2;135;97;60m#[0m[38;2;134;98;60m#[0m[38;2;134;98;61m#[0m[38;2;135;99;60m#[0m[38;2;133;98;58m#[0m[38;2;133;97;58m#[0m[38;2;133;97;58m#[0m");
	$display("[38;2;115;85;49mS[0m[38;2;116;86;49mS[0m[38;2;116;86;49mS[0m[38;2;115;85;49mS[0m[38;2;115;85;49mS[0m[38;2;115;86;49mS[0m[38;2;116;87;50mS[0m[38;2;116;86;50mS[0m[38;2;116;86;50mS[0m[38;2;115;87;50mS[0m[38;2;115;87;50mS[0m[38;2;115;87;50mS[0m[38;2;115;87;50mS[0m[38;2;116;87;50mS[0m[38;2;116;86;50mS[0m[38;2;116;86;50mS[0m[38;2;116;86;50mS[0m[38;2;116;86;50mS[0m[38;2;116;86;50mS[0m[38;2;117;86;48mS[0m[38;2;116;85;48mS[0m[38;2;107;80;48mG[0m[38;2;89;67;41mM[0m[38;2;89;67;44mM[0m[38;2;82;55;29mh[0m[38;2;83;62;41mM[0m[38;2;30;23;11mr[0m[38;2;26;22;14mr[0m[38;2;47;38;28mA[0m[38;2;47;38;31m2[0m[38;2;18;11;8m;[0m[38;2;14;11;9m:[0m[38;2;12;11;8m:[0m[38;2;11;10;7m:[0m[38;2;12;9;7m:[0m[38;2;10;9;8m:[0m[38;2;9;9;7m:[0m[38;2;10;8;6m:[0m[38;2;11;9;10m:[0m[38;2;20;6;7m:[0m[38;2;49;5;4mi[0m[38;2;131;76;65m#[0m[38;2;124;69;58mS[0m[38;2;70;6;8ms[0m[38;2;65;5;9ms[0m[38;2;66;3;8ms[0m[38;2;49;4;7mr[0m[38;2;9;4;2m,[0m[38;2;5;8;7m,[0m[38;2;13;7;7m:[0m[38;2;9;9;6m:[0m[38;2;10;10;8m:[0m[38;2;7;7;5m,[0m[38;2;0;1;0m.[0m[38;2;1;1;1m.[0m[38;2;1;2;1m.[0m[38;2;1;1;2m.[0m[38;2;4;0;0m.[0m[38;2;46;31;28mA[0m[38;2;62;41;34m5[0m[38;2;82;61;47mM[0m[38;2;78;58;43mh[0m[38;2;85;66;53mH[0m[38;2;61;42;32m5[0m[38;2;57;39;31m2[0m[38;2;38;21;18ms[0m[38;2;37;21;19ms[0m[38;2;38;22;20ms[0m[38;2;37;23;20ms[0m[38;2;32;21;20ms[0m[38;2;23;14;13mi[0m[38;2;9;3;2m,[0m[38;2;9;6;5m,[0m[38;2;12;10;9m:[0m[38;2;12;9;8m:[0m[38;2;12;9;9m:[0m[38;2;13;9;9m:[0m[38;2;13;9;10m:[0m[38;2;20;6;5m:[0m[38;2;41;1;2m;[0m[38;2;86;38;34m3[0m[38;2;145;102;87mB[0m[38;2;84;28;23m5[0m[38;2;43;3;4mi[0m[38;2;14;9;6m:[0m[38;2;7;11;10m:[0m[38;2;13;8;10m:[0m[38;2;12;9;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;10;9;7m:[0m[38;2;16;12;11m;[0m[38;2;41;33;26mA[0m[38;2;43;34;27mA[0m[38;2;18;14;12m;[0m[38;2;9;7;6m,[0m[38;2;4;0;0m.[0m[38;2;21;11;7m;[0m[38;2;84;59;42mM[0m[38;2;101;71;43mH[0m[38;2;120;88;53mS[0m[38;2;128;95;59m#[0m[38;2;129;95;61m#[0m[38;2;127;95;58m#[0m[38;2;127;93;57m#[0m[38;2;127;93;57m#[0m[38;2;128;94;58m#[0m[38;2;126;92;57m#[0m[38;2;127;93;56m#[0m[38;2;128;94;57m#[0m[38;2;128;94;56m#[0m[38;2;129;95;57m#[0m[38;2;129;95;57m#[0m[38;2;129;95;58m#[0m[38;2;131;97;60m#[0m[38;2;130;96;59m#[0m[38;2;130;96;59m#[0m[38;2;131;96;59m#[0m[38;2;133;97;59m#[0m[38;2;134;97;60m#[0m[38;2;135;97;60m#[0m[38;2;135;96;59m#[0m[38;2;134;96;59m#[0m[38;2;133;95;58m#[0m[38;2;133;95;57m#[0m[38;2;131;94;55m#[0m[38;2;130;93;55m#[0m[38;2;130;94;56m#[0m");
	$display("[38;2;115;85;49mS[0m[38;2;115;85;49mS[0m[38;2;114;84;48mS[0m[38;2;115;85;49mS[0m[38;2;115;85;49mS[0m[38;2;114;86;49mS[0m[38;2;115;87;50mS[0m[38;2;114;86;49mS[0m[38;2;114;86;49mS[0m[38;2;114;86;49mS[0m[38;2;115;87;50mS[0m[38;2;115;87;50mS[0m[38;2;114;86;49mS[0m[38;2;114;86;49mS[0m[38;2;115;85;49mS[0m[38;2;114;84;48mS[0m[38;2;114;84;48mS[0m[38;2;114;84;48mS[0m[38;2;114;84;48mS[0m[38;2;114;84;48mS[0m[38;2;114;84;48mS[0m[38;2;109;81;50mG[0m[38;2;93;69;41mH[0m[38;2;84;61;36mh[0m[38;2;81;56;27mh[0m[38;2;94;73;47mH[0m[38;2;33;23;12mr[0m[38;2;23;18;14mi[0m[38;2;55;44;32m5[0m[38;2;43;34;24mA[0m[38;2;15;9;8m:[0m[38;2;11;8;8m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;9;9;7m:[0m[38;2;16;5;9m:[0m[38;2;35;2;6m;[0m[38;2;83;36;30m3[0m[38;2;151;100;85mB[0m[38;2;82;21;17m2[0m[38;2;71;4;9ms[0m[38;2;69;2;5ms[0m[38;2;66;2;5ms[0m[38;2;52;3;5mr[0m[38;2;16;2;3m,[0m[38;2;6;6;7m,[0m[38;2;15;10;9m:[0m[38;2;19;15;15mi[0m[38;2;18;15;13m;[0m[38;2;14;14;10m;[0m[38;2;7;6;3m,[0m[38;2;5;2;3m.[0m[38;2;1;1;3m.[0m[38;2;1;1;1m.[0m[38;2;53;39;31m2[0m[38;2;128;105;86m9[0m[38;2;100;81;61mG[0m[38;2;105;86;67mS[0m[38;2;108;85;68mS[0m[38;2;110;85;67mS[0m[38;2;132;108;83m9[0m[38;2;146;119;94mB[0m[38;2;81;57;45mM[0m[38;2;34;18;15mr[0m[38;2;30;17;16mr[0m[38;2;20;14;11m;[0m[38;2;8;7;4m,[0m[38;2;6;5;2m,[0m[38;2;9;7;6m,[0m[38;2;11;9;8m:[0m[38;2;11;10;9m:[0m[38;2;12;10;8m:[0m[38;2;11;10;8m:[0m[38;2;10;10;8m:[0m[38;2;7;8;6m,[0m[38;2;15;5;3m:[0m[38;2;42;3;4mi[0m[38;2;51;0;0mi[0m[38;2;106;60;51mH[0m[38;2;141;96;79m9[0m[38;2;62;13;11mX[0m[38;2;30;5;3m;[0m[38;2;10;9;5m:[0m[38;2;10;10;7m:[0m[38;2;12;9;7m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;10;9;7m:[0m[38;2;15;11;8m:[0m[38;2;46;32;24mA[0m[38;2;54;41;30m2[0m[38;2;24;19;12mi[0m[38;2;6;5;4m,[0m[38;2;3;0;1m.[0m[38;2;35;21;16mr[0m[38;2;85;59;41mM[0m[38;2;99;69;42mH[0m[38;2;116;84;54mS[0m[38;2;124;91;57m#[0m[38;2;125;93;57m#[0m[38;2;123;92;56m#[0m[38;2;124;90;55mS[0m[38;2;124;90;55mS[0m[38;2;124;90;55mS[0m[38;2;124;90;55mS[0m[38;2;125;91;56m#[0m[38;2;125;91;56m#[0m[38;2;125;91;55m#[0m[38;2;125;91;54m#[0m[38;2;126;92;55m#[0m[38;2;126;92;55m#[0m[38;2;127;93;56m#[0m[38;2;127;93;56m#[0m[38;2;127;93;56m#[0m[38;2;127;93;56m#[0m[38;2;129;93;57m#[0m[38;2;129;94;56m#[0m[38;2;129;94;56m#[0m[38;2;129;93;56m#[0m[38;2;129;93;56m#[0m[38;2;129;93;56m#[0m[38;2;129;93;56m#[0m[38;2;128;92;55m#[0m[38;2;127;91;54m#[0m[38;2;127;92;54m#[0m");
	$display("[38;2;114;84;48mS[0m[38;2;114;84;48mS[0m[38;2;114;84;48mS[0m[38;2;114;84;48mS[0m[38;2;114;85;48mS[0m[38;2;114;86;48mS[0m[38;2;114;86;49mS[0m[38;2;114;86;49mS[0m[38;2;114;86;49mS[0m[38;2;114;85;49mS[0m[38;2;115;86;49mS[0m[38;2;114;85;49mS[0m[38;2;113;84;48mS[0m[38;2;113;84;48mS[0m[38;2;113;83;47mG[0m[38;2;113;83;47mG[0m[38;2;113;83;47mG[0m[38;2;113;83;47mG[0m[38;2;113;83;47mG[0m[38;2;113;83;47mG[0m[38;2;113;83;48mG[0m[38;2;110;83;51mG[0m[38;2;95;71;43mH[0m[38;2;79;58;32mh[0m[38;2;88;61;29mh[0m[38;2;107;80;50mG[0m[38;2;54;40;26m2[0m[38;2;18;12;10m;[0m[38;2;57;47;37m5[0m[38;2;57;51;38m5[0m[38;2;19;16;11m;[0m[38;2;9;8;6m:[0m[38;2;9;9;7m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;12;8;8m:[0m[38;2;23;2;3m:[0m[38;2;47;3;3mi[0m[38;2;126;80;71m#[0m[38;2;114;66;56mG[0m[38;2;61;1;1mr[0m[38;2;62;2;5mr[0m[38;2;61;1;2mr[0m[38;2;60;0;5mr[0m[38;2;54;1;5mr[0m[38;2;38;2;8mi[0m[38;2;17;2;4m:[0m[38;2;12;7;5m:[0m[38;2;14;10;10m:[0m[38;2;15;12;9m;[0m[38;2;14;13;8m;[0m[38;2;14;13;8m;[0m[38;2;14;11;10m;[0m[38;2;11;8;9m:[0m[38;2;12;7;5m:[0m[38;2;87;72;61mH[0m[38;2;84;69;52mH[0m[38;2;42;39;24mA[0m[38;2;40;49;32m2[0m[38;2;38;43;23mA[0m[38;2;86;67;49mH[0m[38;2;149;120;98mB[0m[38;2;126;104;82m9[0m[38;2;64;51;41m3[0m[38;2;20;16;13mi[0m[38;2;17;13;10m;[0m[38;2;12;9;5m:[0m[38;2;12;11;7m:[0m[38;2;14;13;10m;[0m[38;2;16;15;13m;[0m[38;2;17;15;13m;[0m[38;2;21;19;18mi[0m[38;2;23;21;20mr[0m[38;2;23;21;18mr[0m[38;2;22;16;14mi[0m[38;2;19;6;6m:[0m[38;2;31;2;4m;[0m[38;2;49;3;8mr[0m[38;2;56;0;3mi[0m[38;2;60;6;3mr[0m[38;2;133;91;78m9[0m[38;2;114;65;56mG[0m[38;2;49;2;2mi[0m[38;2;24;5;5m:[0m[38;2;9;10;7m:[0m[38;2;10;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;11;10;8m:[0m[38;2;10;9;7m:[0m[38;2;26;23;16mr[0m[38;2;67;55;39m3[0m[38;2;60;48;32m5[0m[38;2;19;14;7m;[0m[38;2;4;3;2m.[0m[38;2;5;1;2m.[0m[38;2;46;33;24mA[0m[38;2;82;58;36mh[0m[38;2;96;67;37mM[0m[38;2;112;80;48mG[0m[38;2;122;88;54mS[0m[38;2;123;90;56mS[0m[38;2;120;88;55mS[0m[38;2;122;87;53mS[0m[38;2;122;87;53mS[0m[38;2;122;87;53mS[0m[38;2;121;86;53mS[0m[38;2;121;87;52mS[0m[38;2;122;88;53mS[0m[38;2;122;88;52mS[0m[38;2;123;88;51mS[0m[38;2;123;89;52mS[0m[38;2;124;89;53mS[0m[38;2;126;90;54m#[0m[38;2;125;90;53mS[0m[38;2;126;90;54m#[0m[38;2;126;91;54m#[0m[38;2;126;91;54m#[0m[38;2;126;91;54m#[0m[38;2;126;92;54m#[0m[38;2;126;92;54m#[0m[38;2;126;92;54m#[0m[38;2;126;91;54m#[0m[38;2;126;91;54m#[0m[38;2;125;90;53mS[0m[38;2;124;89;52mS[0m[38;2;125;89;52mS[0m");
	$display("[38;2;113;83;47mG[0m[38;2;113;83;47mG[0m[38;2;113;83;47mG[0m[38;2;113;83;47mG[0m[38;2;113;83;47mG[0m[38;2;113;83;46mG[0m[38;2;112;84;47mG[0m[38;2;111;84;48mG[0m[38;2;112;83;48mG[0m[38;2;112;83;47mG[0m[38;2;112;84;47mG[0m[38;2;112;84;47mG[0m[38;2;112;84;47mG[0m[38;2;112;84;47mG[0m[38;2;112;83;47mG[0m[38;2;111;82;46mG[0m[38;2;111;82;46mG[0m[38;2;111;82;46mG[0m[38;2;112;82;46mG[0m[38;2;112;82;46mG[0m[38;2;111;82;49mG[0m[38;2;107;82;51mG[0m[38;2;95;72;42mH[0m[38;2;79;59;29mh[0m[38;2;90;65;37mM[0m[38;2;108;79;49mG[0m[38;2;83;64;43mM[0m[38;2;17;10;6m:[0m[38;2;30;23;20ms[0m[38;2;31;26;19ms[0m[38;2;13;11;5m:[0m[38;2;9;8;4m,[0m[38;2;9;8;5m,[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;14;7;7m:[0m[38;2;30;2;1m:[0m[38;2;64;20;17mA[0m[38;2;143;98;88m9[0m[38;2;78;29;23m5[0m[38;2;55;0;2mi[0m[38;2;56;0;4mr[0m[38;2;54;1;3mi[0m[38;2;51;1;4mi[0m[38;2;49;1;1mi[0m[38;2;48;2;4mi[0m[38;2;40;2;4m;[0m[38;2;20;2;1m:[0m[38;2;6;5;3m,[0m[38;2;5;7;4m,[0m[38;2;7;8;6m,[0m[38;2;12;10;10m:[0m[38;2;14;10;9m:[0m[38;2;15;9;9m:[0m[38;2;14;10;9m:[0m[38;2;36;29;24mX[0m[38;2;46;40;28mA[0m[38;2;31;34;24mX[0m[38;2;24;34;19ms[0m[38;2;40;46;27mA[0m[38;2;69;56;41mh[0m[38;2;77;60;49mM[0m[38;2;39;30;24mX[0m[38;2;7;3;3m,[0m[38;2;9;10;9m:[0m[38;2;11;10;8m:[0m[38;2;14;11;8m:[0m[38;2;17;13;10m;[0m[38;2;15;11;8m:[0m[38;2;13;9;7m:[0m[38;2;12;8;7m:[0m[38;2;12;9;7m:[0m[38;2;12;8;6m:[0m[38;2;18;3;3m:[0m[38;2;31;1;3m;[0m[38;2;44;3;5mi[0m[38;2;49;2;4mi[0m[38;2;53;1;4mi[0m[38;2;56;0;6mr[0m[38;2;53;0;0mi[0m[38;2;88;39;36m3[0m[38;2;145;103;88mB[0m[38;2;68;19;16mA[0m[38;2;31;2;5m;[0m[38;2;11;7;8m:[0m[38;2;9;9;9m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;10;9;7m:[0m[38;2;9;8;7m:[0m[38;2;10;9;6m:[0m[38;2;10;9;5m:[0m[38;2;10;9;5m:[0m[38;2;10;8;5m:[0m[38;2;19;15;11m;[0m[38;2;41;35;25mA[0m[38;2;30;25;17mr[0m[38;2;10;6;6m,[0m[38;2;4;1;2m.[0m[38;2;15;10;6m:[0m[38;2;58;42;26m2[0m[38;2;79;59;31mh[0m[38;2;91;66;36mM[0m[38;2;106;77;46mG[0m[38;2;114;84;51mS[0m[38;2;115;85;52mS[0m[38;2;112;82;52mS[0m[38;2;113;81;51mS[0m[38;2;112;82;51mS[0m[38;2;111;82;51mG[0m[38;2;111;81;50mG[0m[38;2;111;81;48mG[0m[38;2;113;82;49mG[0m[38;2;115;83;49mS[0m[38;2;114;83;49mS[0m[38;2;113;83;49mS[0m[38;2;114;83;48mS[0m[38;2;116;84;50mS[0m[38;2;116;85;50mS[0m[38;2;115;84;49mS[0m[38;2;115;84;49mS[0m[38;2;115;84;49mS[0m[38;2;115;84;49mS[0m[38;2;115;84;49mS[0m[38;2;115;84;49mS[0m[38;2;115;83;49mS[0m[38;2;115;84;49mS[0m[38;2;115;83;49mS[0m[38;2;115;83;48mS[0m[38;2;115;82;48mS[0m[38;2;114;82;48mG[0m");
	$display("\033[0;32m \033[5m    //   ) )     // | |     //   ) )     //   ) )\033[m");
    $display("\033[0;32m \033[5m   //___/ /     //__| |    ((           ((\033[m");
    $display("\033[0;32m \033[5m  / ____ /     / ___  |      \\           \\\033[m");
    $display("\033[0;32m \033[5m //           //    | |        ) )          ) )\033[m");
    $display("\033[0;32m \033[5m//           //     | | ((___ / /    ((___ / /\033[m");
	$display("**************************************************");
	$display("                  Congratulations!                ");
	$display("              execution cycles = %7d", total_latency);
	$display("              clock period = %4fns", CYCLE);
	$display("**************************************************");
end endtask

endmodule